
//Verilog file of module CPU


`timescale 1 ns / 1ns

module CPU_net(
inst,
CPU_wire_75,CPU_wire_78,CPU_wire_86,CPU_wire_88,CPU_wire_2,CPU_wire_4,CPU_wire_92,CPU_wire_7,
CPU_wire_126,CPU_wire_142,CPU_wire_158,CPU_wire_174,CPU_wire_190,CPU_wire_206,CPU_wire_222,CPU_wire_238,CPU_wire_116,
CPU_wire_132,CPU_wire_148,CPU_wire_164,CPU_wire_180,CPU_wire_196, CPU_wire_212,CPU_wire_228,CPU_wire_123,CPU_wire_139,
CPU_wire_155,CPU_wire_171,CPU_wire_187,CPU_wire_203,CPU_wire_219,CPU_wire_235,CPU_wire_112, CPU_wire_128,CPU_wire_144,
CPU_wire_160,CPU_wire_176,CPU_wire_192,CPU_wire_208,CPU_wire_224,CPU_wire_10,CPU_wire_12,CPU_wire_14,CPU_wire_16,CPU_wire_18,
CPU_wire_20,CPU_wire_22,CPU_wire_24,CPU_wire_58,CPU_wire_61,CPU_wire_63,CPU_wire_65,CPU_wire_67,CPU_wire_69,CPU_wire_71,
CPU_wire_73,
address,
out_data,
store,
CPU_wire_83,CPU_wire_84,CPU_wire_85,CPU_wire_87,CPU_wire_89,CPU_wire_90,CPU_wire_91,CPU_wire_93,
CPU_wire_337,CPU_wire_338,CPU_wire_339,CPU_wire_340,CPU_wire_341,CPU_wire_342,CPU_wire_343,CPU_wire_344,CPU_wire_346,CPU_wire_347,CPU_wire_348,CPU_wire_349,
CPU_wire_350,CPU_wire_351,CPU_wire_352,CPU_wire_353,CPU_wire_355,CPU_wire_356,CPU_wire_357,CPU_wire_358,CPU_wire_359,CPU_wire_360,CPU_wire_361,CPU_wire_362,
CPU_wire_364,CPU_wire_365,CPU_wire_366,CPU_wire_367,CPU_wire_368,CPU_wire_369,CPU_wire_370,CPU_wire_371,CPU_wire_501,CPU_wire_503,CPU_wire_505,CPU_wire_507,
CPU_wire_509,CPU_wire_511,CPU_wire_513,CPU_wire_515,CPU_wire_619,CPU_wire_622,CPU_wire_625,CPU_wire_628,CPU_wire_631,CPU_wire_634,CPU_wire_637,CPU_wire_640
);
	
	input CPU_wire_75,CPU_wire_78,CPU_wire_86,CPU_wire_88,CPU_wire_2,CPU_wire_4,CPU_wire_92,CPU_wire_7,
CPU_wire_126,CPU_wire_142,CPU_wire_158,CPU_wire_174,CPU_wire_190,CPU_wire_206,CPU_wire_222,CPU_wire_238,CPU_wire_116,
CPU_wire_132,CPU_wire_148,CPU_wire_164,CPU_wire_180,CPU_wire_196, CPU_wire_212,CPU_wire_228,CPU_wire_123,CPU_wire_139,
CPU_wire_155,CPU_wire_171,CPU_wire_187,CPU_wire_203,CPU_wire_219,CPU_wire_235,CPU_wire_112, CPU_wire_128,CPU_wire_144,
CPU_wire_160,CPU_wire_176,CPU_wire_192,CPU_wire_208,CPU_wire_224,CPU_wire_10,CPU_wire_12,CPU_wire_14,CPU_wire_16,CPU_wire_18,
CPU_wire_20,CPU_wire_22,CPU_wire_24,CPU_wire_58,CPU_wire_61,CPU_wire_63,CPU_wire_65,CPU_wire_67,CPU_wire_69,CPU_wire_71,CPU_wire_73;

input [0:7]inst;
output [0:7]address;
output [0:7]out_data;
    output store;
	output CPU_wire_83,CPU_wire_84,CPU_wire_85,CPU_wire_87,CPU_wire_89,CPU_wire_90,CPU_wire_91,CPU_wire_93,
CPU_wire_337,CPU_wire_338,CPU_wire_339,CPU_wire_340,CPU_wire_341,CPU_wire_342,CPU_wire_343,CPU_wire_344,CPU_wire_346,CPU_wire_347,CPU_wire_348,CPU_wire_349,
CPU_wire_350,CPU_wire_351,CPU_wire_352,CPU_wire_353,CPU_wire_355,CPU_wire_356,CPU_wire_357,CPU_wire_358,CPU_wire_359,CPU_wire_360,CPU_wire_361,CPU_wire_362,
CPU_wire_364,CPU_wire_365,CPU_wire_366,CPU_wire_367,CPU_wire_368,CPU_wire_369,CPU_wire_370,CPU_wire_371,CPU_wire_501,CPU_wire_503,CPU_wire_505,CPU_wire_507,
CPU_wire_509,CPU_wire_511,CPU_wire_513,CPU_wire_515,CPU_wire_619,CPU_wire_622,CPU_wire_625,CPU_wire_628,CPU_wire_631,CPU_wire_634,CPU_wire_637,CPU_wire_640;

wire
CPU_wire_1,
CPU_wire_2,
CPU_wire_3,
CPU_wire_4,
CPU_wire_5,
CPU_wire_6,
CPU_wire_7,
CPU_wire_8,
CPU_wire_9,
CPU_wire_10,
CPU_wire_11,
CPU_wire_12,
CPU_wire_13,
CPU_wire_14,
CPU_wire_15,
CPU_wire_16,
CPU_wire_17,
CPU_wire_18,
CPU_wire_19,
CPU_wire_20,
CPU_wire_21,
CPU_wire_22,
CPU_wire_23,
CPU_wire_24,
CPU_wire_25,
CPU_wire_26,
CPU_wire_27,
CPU_wire_28,
CPU_wire_29,
CPU_wire_30,
CPU_wire_31,
CPU_wire_32,
CPU_wire_33,
CPU_wire_34,
CPU_wire_35,
CPU_wire_36,
CPU_wire_37,
CPU_wire_38,
CPU_wire_39,
CPU_wire_40,
CPU_wire_41,
CPU_wire_42,
CPU_wire_43,
CPU_wire_44,
CPU_wire_45,
CPU_wire_46,
CPU_wire_47,
CPU_wire_48,
CPU_wire_49,
CPU_wire_50,
CPU_wire_51,
CPU_wire_52,
CPU_wire_53,
CPU_wire_54,
CPU_wire_55,
CPU_wire_56,
CPU_wire_57,
CPU_wire_58,
CPU_wire_59,
CPU_wire_60,
CPU_wire_61,
CPU_wire_62,
CPU_wire_63,
CPU_wire_64,
CPU_wire_65,
CPU_wire_66,
CPU_wire_67,
CPU_wire_68,
CPU_wire_69,
CPU_wire_70,
CPU_wire_71,
CPU_wire_72,
CPU_wire_73,
CPU_wire_74,
CPU_wire_75,
CPU_wire_76,
CPU_wire_77,
CPU_wire_78,
CPU_wire_79,
CPU_wire_80,
CPU_wire_81,
CPU_wire_82,
CPU_wire_83,
CPU_wire_84,
CPU_wire_85,
CPU_wire_86,
CPU_wire_87,
CPU_wire_88,
CPU_wire_89,
CPU_wire_90,
CPU_wire_91,
CPU_wire_92,
CPU_wire_93,
CPU_wire_94,
CPU_wire_95,
CPU_wire_96,
CPU_wire_97,
CPU_wire_98,
CPU_wire_99,
CPU_wire_100,
CPU_wire_101,
CPU_wire_102,
CPU_wire_103,
CPU_wire_104,
CPU_wire_105,
CPU_wire_106,
CPU_wire_107,
CPU_wire_108,
CPU_wire_109,
CPU_wire_110,
CPU_wire_111,
CPU_wire_112,
CPU_wire_113,
CPU_wire_114,
CPU_wire_115,
CPU_wire_116,
CPU_wire_117,
CPU_wire_118,
CPU_wire_119,
CPU_wire_120,
CPU_wire_121,
CPU_wire_122,
CPU_wire_123,
CPU_wire_124,
CPU_wire_125,
CPU_wire_126,
CPU_wire_127,
CPU_wire_128,
CPU_wire_129,
CPU_wire_130,
CPU_wire_131,
CPU_wire_132,
CPU_wire_133,
CPU_wire_134,
CPU_wire_135,
CPU_wire_136,
CPU_wire_137,
CPU_wire_138,
CPU_wire_139,
CPU_wire_140,
CPU_wire_141,
CPU_wire_142,
CPU_wire_143,
CPU_wire_144,
CPU_wire_145,
CPU_wire_146,
CPU_wire_147,
CPU_wire_148,
CPU_wire_149,
CPU_wire_150,
CPU_wire_151,
CPU_wire_152,
CPU_wire_153,
CPU_wire_154,
CPU_wire_155,
CPU_wire_156,
CPU_wire_157,
CPU_wire_158,
CPU_wire_159,
CPU_wire_160,
CPU_wire_161,
CPU_wire_162,
CPU_wire_163,
CPU_wire_164,
CPU_wire_165,
CPU_wire_166,
CPU_wire_167,
CPU_wire_168,
CPU_wire_169,
CPU_wire_170,
CPU_wire_171,
CPU_wire_172,
CPU_wire_173,
CPU_wire_174,
CPU_wire_175,
CPU_wire_176,
CPU_wire_177,
CPU_wire_178,
CPU_wire_179,
CPU_wire_180,
CPU_wire_181,
CPU_wire_182,
CPU_wire_183,
CPU_wire_184,
CPU_wire_185,
CPU_wire_186,
CPU_wire_187,
CPU_wire_188,
CPU_wire_189,
CPU_wire_190,
CPU_wire_191,
CPU_wire_192,
CPU_wire_193,
CPU_wire_194,
CPU_wire_195,
CPU_wire_196,
CPU_wire_197,
CPU_wire_198,
CPU_wire_199,
CPU_wire_200,
CPU_wire_201,
CPU_wire_202,
CPU_wire_203,
CPU_wire_204,
CPU_wire_205,
CPU_wire_206,
CPU_wire_207,
CPU_wire_208,
CPU_wire_209,
CPU_wire_210,
CPU_wire_211,
CPU_wire_212,
CPU_wire_213,
CPU_wire_214,
CPU_wire_215,
CPU_wire_216,
CPU_wire_217,
CPU_wire_218,
CPU_wire_219,
CPU_wire_220,
CPU_wire_221,
CPU_wire_222,
CPU_wire_223,
CPU_wire_224,
CPU_wire_225,
CPU_wire_226,
CPU_wire_227,
CPU_wire_228,
CPU_wire_229,
CPU_wire_230,
CPU_wire_231,
CPU_wire_232,
CPU_wire_233,
CPU_wire_234,
CPU_wire_235,
CPU_wire_236,
CPU_wire_237,
CPU_wire_238,
CPU_wire_239,
CPU_wire_240,
CPU_wire_241,
CPU_wire_242,
CPU_wire_243,
CPU_wire_244,
CPU_wire_245,
CPU_wire_246,
CPU_wire_247,
CPU_wire_248,
CPU_wire_249,
CPU_wire_250,
CPU_wire_251,
CPU_wire_252,
CPU_wire_253,
CPU_wire_254,
CPU_wire_255,
CPU_wire_256,
CPU_wire_257,
CPU_wire_258,
CPU_wire_259,
CPU_wire_260,
CPU_wire_261,
CPU_wire_262,
CPU_wire_263,
CPU_wire_264,
CPU_wire_265,
CPU_wire_266,
CPU_wire_267,
CPU_wire_268,
CPU_wire_269,
CPU_wire_270,
CPU_wire_271,
CPU_wire_272,
CPU_wire_273,
CPU_wire_274,
CPU_wire_275,
CPU_wire_276,
CPU_wire_277,
CPU_wire_278,
CPU_wire_279,
CPU_wire_280,
CPU_wire_281,
CPU_wire_282,
CPU_wire_283,
CPU_wire_284,
CPU_wire_285,
CPU_wire_286,
CPU_wire_287,
CPU_wire_288,
CPU_wire_289,
CPU_wire_290,
CPU_wire_291,
CPU_wire_292,
CPU_wire_293,
CPU_wire_294,
CPU_wire_295,
CPU_wire_296,
CPU_wire_297,
CPU_wire_298,
CPU_wire_299,
CPU_wire_300,
CPU_wire_301,
CPU_wire_302,
CPU_wire_303,
CPU_wire_304,
CPU_wire_305,
CPU_wire_306,
CPU_wire_307,
CPU_wire_308,
CPU_wire_309,
CPU_wire_310,
CPU_wire_311,
CPU_wire_312,
CPU_wire_313,
CPU_wire_314,
CPU_wire_315,
CPU_wire_316,
CPU_wire_317,
CPU_wire_318,
CPU_wire_319,
CPU_wire_320,
CPU_wire_321,
CPU_wire_322,
CPU_wire_323,
CPU_wire_324,
CPU_wire_325,
CPU_wire_326,
CPU_wire_327,
CPU_wire_328,
CPU_wire_329,
CPU_wire_330,
CPU_wire_331,
CPU_wire_332,
CPU_wire_333,
CPU_wire_334,
CPU_wire_335,
CPU_wire_336,
CPU_wire_337,
CPU_wire_338,
CPU_wire_339,
CPU_wire_340,
CPU_wire_341,
CPU_wire_342,
CPU_wire_343,
CPU_wire_344,
CPU_wire_345,
CPU_wire_346,
CPU_wire_347,
CPU_wire_348,
CPU_wire_349,
CPU_wire_350,
CPU_wire_351,
CPU_wire_352,
CPU_wire_353,
CPU_wire_354,
CPU_wire_355,
CPU_wire_356,
CPU_wire_357,
CPU_wire_358,
CPU_wire_359,
CPU_wire_360,
CPU_wire_361,
CPU_wire_362,
CPU_wire_363,
CPU_wire_364,
CPU_wire_365,
CPU_wire_366,
CPU_wire_367,
CPU_wire_368,
CPU_wire_369,
CPU_wire_370,
CPU_wire_371,
CPU_wire_372,
CPU_wire_373,
CPU_wire_374,
CPU_wire_375,
CPU_wire_376,
CPU_wire_377,
CPU_wire_378,
CPU_wire_379,
CPU_wire_380,
CPU_wire_381,
CPU_wire_382,
CPU_wire_383,
CPU_wire_384,
CPU_wire_385,
CPU_wire_386,
CPU_wire_387,
CPU_wire_388,
CPU_wire_389,
CPU_wire_390,
CPU_wire_391,
CPU_wire_392,
CPU_wire_393,
CPU_wire_394,
CPU_wire_395,
CPU_wire_396,
CPU_wire_397,
CPU_wire_398,
CPU_wire_399,
CPU_wire_400,
CPU_wire_401,
CPU_wire_402,
CPU_wire_403,
CPU_wire_404,
CPU_wire_405,
CPU_wire_406,
CPU_wire_407,
CPU_wire_408,
CPU_wire_409,
CPU_wire_410,
CPU_wire_411,
CPU_wire_412,
CPU_wire_413,
CPU_wire_414,
CPU_wire_415,
CPU_wire_416,
CPU_wire_417,
CPU_wire_418,
CPU_wire_419,
CPU_wire_420,
CPU_wire_421,
CPU_wire_422,
CPU_wire_423,
CPU_wire_424,
CPU_wire_425,
CPU_wire_426,
CPU_wire_427,
CPU_wire_428,
CPU_wire_429,
CPU_wire_430,
CPU_wire_431,
CPU_wire_432,
CPU_wire_433,
CPU_wire_434,
CPU_wire_435,
CPU_wire_436,
CPU_wire_437,
CPU_wire_438,
CPU_wire_439,
CPU_wire_440,
CPU_wire_441,
CPU_wire_442,
CPU_wire_443,
CPU_wire_444,
CPU_wire_445,
CPU_wire_446,
CPU_wire_447,
CPU_wire_448,
CPU_wire_449,
CPU_wire_450,
CPU_wire_451,
CPU_wire_452,
CPU_wire_453,
CPU_wire_454,
CPU_wire_455,
CPU_wire_456,
CPU_wire_457,
CPU_wire_458,
CPU_wire_459,
CPU_wire_460,
CPU_wire_461,
CPU_wire_462,
CPU_wire_463,
CPU_wire_464,
CPU_wire_465,
CPU_wire_466,
CPU_wire_467,
CPU_wire_468,
CPU_wire_469,
CPU_wire_470,
CPU_wire_471,
CPU_wire_472,
CPU_wire_473,
CPU_wire_474,
CPU_wire_475,
CPU_wire_476,
CPU_wire_477,
CPU_wire_478,
CPU_wire_479,
CPU_wire_480,
CPU_wire_481,
CPU_wire_482,
CPU_wire_483,
CPU_wire_484,
CPU_wire_485,
CPU_wire_486,
CPU_wire_487,
CPU_wire_488,
CPU_wire_489,
CPU_wire_490,
CPU_wire_491,
CPU_wire_492,
CPU_wire_493,
CPU_wire_494,
CPU_wire_495,
CPU_wire_496,
CPU_wire_497,
CPU_wire_498,
CPU_wire_499,
CPU_wire_500,
CPU_wire_501,
CPU_wire_502,
CPU_wire_503,
CPU_wire_504,
CPU_wire_505,
CPU_wire_506,
CPU_wire_507,
CPU_wire_508,
CPU_wire_509,
CPU_wire_510,
CPU_wire_511,
CPU_wire_512,
CPU_wire_513,
CPU_wire_514,
CPU_wire_515,
CPU_wire_516,
CPU_wire_517,
CPU_wire_518,
CPU_wire_519,
CPU_wire_520,
CPU_wire_521,
CPU_wire_522,
CPU_wire_523,
CPU_wire_524,
CPU_wire_525,
CPU_wire_526,
CPU_wire_527,
CPU_wire_528,
CPU_wire_529,
CPU_wire_530,
CPU_wire_531,
CPU_wire_532,
CPU_wire_533,
CPU_wire_534,
CPU_wire_535,
CPU_wire_536,
CPU_wire_537,
CPU_wire_538,
CPU_wire_539,
CPU_wire_540,
CPU_wire_541,
CPU_wire_542,
CPU_wire_543,
CPU_wire_544,
CPU_wire_545,
CPU_wire_546,
CPU_wire_547,
CPU_wire_548,
CPU_wire_549,
CPU_wire_550,
CPU_wire_551,
CPU_wire_552,
CPU_wire_553,
CPU_wire_554,
CPU_wire_555,
CPU_wire_556,
CPU_wire_557,
CPU_wire_558,
CPU_wire_559,
CPU_wire_560,
CPU_wire_561,
CPU_wire_562,
CPU_wire_563,
CPU_wire_564,
CPU_wire_565,
CPU_wire_566,
CPU_wire_567,
CPU_wire_568,
CPU_wire_569,
CPU_wire_570,
CPU_wire_571,
CPU_wire_572,
CPU_wire_573,
CPU_wire_574,
CPU_wire_575,
CPU_wire_576,
CPU_wire_577,
CPU_wire_578,
CPU_wire_579,
CPU_wire_580,
CPU_wire_581,
CPU_wire_582,
CPU_wire_583,
CPU_wire_584,
CPU_wire_585,
CPU_wire_586,
CPU_wire_587,
CPU_wire_588,
CPU_wire_589,
CPU_wire_590,
CPU_wire_591,
CPU_wire_592,
CPU_wire_593,
CPU_wire_594,
CPU_wire_595,
CPU_wire_596,
CPU_wire_597,
CPU_wire_598,
CPU_wire_599,
CPU_wire_600,
CPU_wire_601,
CPU_wire_602,
CPU_wire_603,
CPU_wire_604,
CPU_wire_605,
CPU_wire_606,
CPU_wire_607,
CPU_wire_608,
CPU_wire_609,
CPU_wire_610,
CPU_wire_611,
CPU_wire_612,
CPU_wire_613,
CPU_wire_614,
CPU_wire_615,
CPU_wire_616,
CPU_wire_617,
CPU_wire_618,
CPU_wire_619,
CPU_wire_620,
CPU_wire_621,
CPU_wire_622,
CPU_wire_623,
CPU_wire_624,
CPU_wire_625,
CPU_wire_626,
CPU_wire_627,
CPU_wire_628,
CPU_wire_629,
CPU_wire_630,
CPU_wire_631,
CPU_wire_632,
CPU_wire_633,
CPU_wire_634,
CPU_wire_635,
CPU_wire_636,
CPU_wire_637,
CPU_wire_638,
CPU_wire_639,
CPU_wire_640,
CPU_wire_641,
CPU_wire_642,
CPU_wire_643,
CPU_wire_644,
CPU_wire_645,
CPU_wire_646,
CPU_wire_647,
CPU_wire_648,
CPU_wire_649,
CPU_wire_650,
CPU_wire_651,
CPU_wire_652,
CPU_wire_653,
CPU_wire_654,
CPU_wire_655,
CPU_wire_656,
CPU_wire_657,
CPU_wire_658,
CPU_wire_659,
CPU_wire_660,
CPU_wire_661,
CPU_wire_662,
CPU_wire_663,
CPU_wire_664,
CPU_wire_665,
CPU_wire_666,
CPU_wire_667,
CPU_wire_668,
CPU_wire_669,
CPU_wire_670,
CPU_wire_671,
CPU_wire_672,
CPU_wire_673,
CPU_wire_674,
CPU_wire_675,
CPU_wire_676,
CPU_wire_677,
CPU_wire_678,
CPU_wire_679,
CPU_wire_680,
CPU_wire_681,
CPU_wire_682,
CPU_wire_683,
CPU_wire_684,
CPU_wire_685,
CPU_wire_686,
CPU_wire_687,
CPU_wire_688,
CPU_wire_689,
CPU_wire_690,
CPU_wire_691,
CPU_wire_692,
CPU_wire_693,
CPU_wire_694,
CPU_wire_695,
CPU_wire_696,
CPU_wire_697,
CPU_wire_698,
CPU_wire_699,
CPU_wire_700,
CPU_wire_701,
CPU_wire_702,
CPU_wire_703,
CPU_wire_704,
CPU_wire_705,
CPU_wire_706,
CPU_wire_707,
CPU_wire_708,
CPU_wire_709,
CPU_wire_710,
CPU_wire_711,
CPU_wire_712,
CPU_wire_713,
CPU_wire_714,
CPU_wire_715,
CPU_wire_716,
CPU_wire_717,
CPU_wire_718,
CPU_wire_719,
CPU_wire_720,
CPU_wire_721,
CPU_wire_722,
CPU_wire_723,
CPU_wire_724,
CPU_wire_725,
CPU_wire_726,
CPU_wire_727,
CPU_wire_728,
CPU_wire_729,
CPU_wire_730,
CPU_wire_731,
CPU_wire_732,
CPU_wire_733,
CPU_wire_734,
CPU_wire_735,
CPU_wire_736,
CPU_wire_737,
CPU_wire_738,
CPU_wire_739,
CPU_wire_740,
CPU_wire_741,
CPU_wire_742,
CPU_wire_743,
CPU_wire_744,
CPU_wire_745,
CPU_wire_746,
CPU_wire_6_0,
CPU_wire_6_1,
CPU_wire_6_2,
CPU_wire_6_3,
CPU_wire_6_4,
CPU_wire_6_5,
CPU_wire_6_6,
CPU_wire_6_7,
CPU_wire_6_8,
CPU_wire_6_9,
CPU_wire_6_10,
CPU_wire_6_11,
CPU_wire_6_12,
CPU_wire_6_13,
CPU_wire_6_14,
CPU_wire_6_15,
CPU_wire_6_16,
CPU_wire_6_17,
CPU_wire_6_18,
CPU_wire_6_19,
CPU_wire_6_20,
CPU_wire_6_21,
CPU_wire_6_22,
CPU_wire_6_23,
CPU_wire_6_24,
CPU_wire_6_25,
CPU_wire_6_26,
CPU_wire_6_27,
CPU_wire_6_28,
CPU_wire_6_29,
CPU_wire_6_30,
CPU_wire_6_31,
CPU_wire_8_0,
CPU_wire_8_1,
CPU_wire_8_2,
CPU_wire_8_3,
CPU_wire_8_4,
CPU_wire_8_5,
CPU_wire_8_6,
CPU_wire_8_7,
CPU_wire_8_8,
CPU_wire_8_9,
CPU_wire_8_10,
CPU_wire_8_11,
CPU_wire_8_12,
CPU_wire_8_13,
CPU_wire_8_14,
CPU_wire_8_15,
CPU_wire_8_16,
CPU_wire_8_17,
CPU_wire_8_18,
CPU_wire_8_19,
CPU_wire_8_20,
CPU_wire_8_21,
CPU_wire_8_22,
CPU_wire_8_23,
CPU_wire_8_24,
CPU_wire_8_25,
CPU_wire_8_26,
CPU_wire_8_27,
CPU_wire_8_28,
CPU_wire_8_29,
CPU_wire_8_30,
CPU_wire_8_31,
CPU_wire_8_32,
CPU_wire_8_33,
CPU_wire_8_34,
CPU_wire_8_35,
CPU_wire_49_0,
CPU_wire_49_1,
CPU_wire_50_0,
CPU_wire_50_1,
CPU_wire_51_0,
CPU_wire_51_1,
CPU_wire_52_0,
CPU_wire_52_1,
CPU_wire_53_0,
CPU_wire_53_1,
CPU_wire_54_0,
CPU_wire_54_1,
CPU_wire_55_0,
CPU_wire_55_1,
CPU_wire_56_0,
CPU_wire_56_1,
CPU_wire_62_0,
CPU_wire_62_1,
CPU_wire_62_2,
CPU_wire_62_3,
CPU_wire_64_0,
CPU_wire_64_1,
CPU_wire_64_2,
CPU_wire_64_3,
CPU_wire_66_0,
CPU_wire_66_1,
CPU_wire_66_2,
CPU_wire_66_3,
CPU_wire_68_0,
CPU_wire_68_1,
CPU_wire_68_2,
CPU_wire_68_3,
CPU_wire_70_0,
CPU_wire_70_1,
CPU_wire_70_2,
CPU_wire_70_3,
CPU_wire_72_0,
CPU_wire_72_1,
CPU_wire_72_2,
CPU_wire_72_3,
CPU_wire_80_0,
CPU_wire_80_1,
CPU_wire_80_2,
CPU_wire_80_3,
CPU_wire_81_0,
CPU_wire_81_1,
CPU_wire_81_2,
CPU_wire_81_3,
CPU_wire_75_0,
CPU_wire_75_1,
CPU_wire_75_2,
CPU_wire_75_3,
CPU_wire_75_4,
CPU_wire_75_5,
CPU_wire_75_6,
CPU_wire_75_7,
CPU_wire_75_8,
CPU_wire_75_9,
CPU_wire_75_10,
CPU_wire_75_11,
CPU_wire_75_12,
CPU_wire_75_13,
CPU_wire_75_14,
CPU_wire_75_15,
CPU_wire_75_16,
CPU_wire_75_17,
CPU_wire_75_18,
CPU_wire_78_0,
CPU_wire_78_1,
CPU_wire_78_2,
CPU_wire_78_3,
CPU_wire_78_4,
CPU_wire_78_5,
CPU_wire_78_6,
CPU_wire_78_7,
CPU_wire_78_8,
CPU_wire_78_9,
CPU_wire_78_10,
CPU_wire_78_11,
CPU_wire_78_12,
CPU_wire_78_13,
CPU_wire_78_14,
CPU_wire_78_15,
CPU_wire_78_16,
CPU_wire_78_17,
CPU_wire_78_18,
CPU_wire_78_19,
CPU_wire_78_20,
CPU_wire_78_21,
CPU_wire_78_22,
CPU_wire_78_23,
CPU_wire_78_24,
CPU_wire_78_25,
CPU_wire_78_26,
CPU_wire_78_27,
CPU_wire_78_28,
CPU_wire_78_29,
CPU_wire_78_30,
CPU_wire_78_31,
CPU_wire_78_32,
CPU_wire_78_33,
CPU_wire_78_34,
CPU_wire_78_35,
CPU_wire_86_0,
CPU_wire_86_1,
CPU_wire_86_2,
CPU_wire_86_3,
CPU_wire_86_4,
CPU_wire_86_5,
CPU_wire_86_6,
CPU_wire_86_7,
CPU_wire_86_8,
CPU_wire_86_9,
CPU_wire_86_10,
CPU_wire_86_11,
CPU_wire_86_12,
CPU_wire_86_13,
CPU_wire_86_14,
CPU_wire_86_15,
CPU_wire_86_16,
CPU_wire_86_17,
CPU_wire_86_18,
CPU_wire_86_19,
CPU_wire_86_20,
CPU_wire_86_21,
CPU_wire_86_22,
CPU_wire_86_23,
CPU_wire_86_24,
CPU_wire_86_25,
CPU_wire_86_26,
CPU_wire_86_27,
CPU_wire_86_28,
CPU_wire_86_29,
CPU_wire_86_30,
CPU_wire_86_31,
CPU_wire_86_32,
CPU_wire_86_33,
CPU_wire_86_34,
CPU_wire_86_35,
CPU_wire_86_36,
CPU_wire_86_37,
CPU_wire_86_38,
CPU_wire_86_39,
CPU_wire_86_40,
CPU_wire_86_41,
CPU_wire_86_42,
CPU_wire_86_43,
CPU_wire_86_44,
CPU_wire_86_45,
CPU_wire_86_46,
CPU_wire_86_47,
CPU_wire_86_48,
CPU_wire_86_49,
CPU_wire_86_50,
CPU_wire_86_51,
CPU_wire_86_52,
CPU_wire_86_53,
CPU_wire_86_54,
CPU_wire_88_0,
CPU_wire_88_1,
CPU_wire_88_2,
CPU_wire_88_3,
CPU_wire_88_4,
CPU_wire_88_5,
CPU_wire_88_6,
CPU_wire_88_7,
CPU_wire_88_8,
CPU_wire_88_9,
CPU_wire_88_10,
CPU_wire_88_11,
CPU_wire_88_12,
CPU_wire_88_13,
CPU_wire_88_14,
CPU_wire_88_15,
CPU_wire_88_16,
CPU_wire_88_17,
CPU_wire_88_18,
CPU_wire_88_19,
CPU_wire_88_20,
CPU_wire_88_21,
CPU_wire_88_22,
CPU_wire_88_23,
CPU_wire_88_24,
CPU_wire_88_25,
CPU_wire_88_26,
CPU_wire_88_27,
CPU_wire_88_28,
CPU_wire_88_29,
CPU_wire_88_30,
CPU_wire_88_31,
CPU_wire_88_32,
CPU_wire_88_33,
CPU_wire_88_34,
CPU_wire_88_35,
CPU_wire_88_36,
CPU_wire_88_37,
CPU_wire_88_38,
CPU_wire_88_39,
CPU_wire_88_40,
CPU_wire_88_41,
CPU_wire_88_42,
CPU_wire_88_43,
CPU_wire_88_44,
CPU_wire_88_45,
CPU_wire_88_46,
CPU_wire_88_47,
CPU_wire_88_48,
CPU_wire_88_49,
CPU_wire_88_50,
CPU_wire_88_51,
CPU_wire_88_52,
CPU_wire_88_53,
CPU_wire_88_54,
CPU_wire_88_55,
CPU_wire_88_56,
CPU_wire_88_57,
CPU_wire_88_58,
CPU_wire_88_59,
CPU_wire_88_60,
CPU_wire_88_61,
CPU_wire_88_62,
CPU_wire_88_63,
CPU_wire_88_64,
CPU_wire_88_65,
CPU_wire_88_66,
CPU_wire_88_67,
CPU_wire_88_68,
CPU_wire_88_69,
CPU_wire_88_70,
CPU_wire_2_0,
CPU_wire_2_1,
CPU_wire_2_2,
CPU_wire_2_3,
CPU_wire_2_4,
CPU_wire_2_5,
CPU_wire_2_6,
CPU_wire_2_7,
CPU_wire_2_8,
CPU_wire_2_9,
CPU_wire_2_10,
CPU_wire_2_11,
CPU_wire_4_0,
CPU_wire_4_1,
CPU_wire_4_2,
CPU_wire_4_3,
CPU_wire_4_4,
CPU_wire_4_5,
CPU_wire_4_6,
CPU_wire_4_7,
CPU_wire_4_8,
CPU_wire_4_9,
CPU_wire_4_10,
CPU_wire_4_11,
CPU_wire_4_12,
CPU_wire_7_0,
CPU_wire_7_1,
CPU_wire_7_2,
CPU_wire_7_3,
CPU_wire_7_4,
CPU_wire_7_5,
CPU_wire_7_6,
CPU_wire_7_7,
CPU_wire_7_8,
CPU_wire_7_9,
CPU_wire_7_10,
CPU_wire_7_11,
CPU_wire_7_12,
CPU_wire_7_13,
CPU_wire_7_14,
CPU_wire_7_15,
CPU_wire_7_16,
CPU_wire_7_17,
CPU_wire_120_0,
CPU_wire_120_1,
CPU_wire_120_2,
CPU_wire_136_0,
CPU_wire_136_1,
CPU_wire_136_2,
CPU_wire_136_3,
CPU_wire_136_4,
CPU_wire_136_5,
CPU_wire_136_6,
CPU_wire_152_0,
CPU_wire_152_1,
CPU_wire_152_2,
CPU_wire_152_3,
CPU_wire_152_4,
CPU_wire_168_0,
CPU_wire_168_1,
CPU_wire_168_2,
CPU_wire_168_3,
CPU_wire_168_4,
CPU_wire_184_0,
CPU_wire_184_1,
CPU_wire_184_2,
CPU_wire_184_3,
CPU_wire_184_4,
CPU_wire_200_0,
CPU_wire_200_1,
CPU_wire_200_2,
CPU_wire_200_3,
CPU_wire_200_4,
CPU_wire_216_0,
CPU_wire_216_1,
CPU_wire_216_2,
CPU_wire_216_3,
CPU_wire_216_4,
CPU_wire_232_0,
CPU_wire_232_1,
CPU_wire_232_2,
CPU_wire_232_3,
CPU_wire_232_4,
CPU_wire_246_0,
CPU_wire_246_1,
CPU_wire_258_0,
CPU_wire_258_1,
CPU_wire_258_2,
CPU_wire_258_3,
CPU_wire_258_4,
CPU_wire_258_5,
CPU_wire_270_0,
CPU_wire_270_1,
CPU_wire_270_2,
CPU_wire_270_3,
CPU_wire_270_4,
CPU_wire_270_5,
CPU_wire_282_0,
CPU_wire_282_1,
CPU_wire_282_2,
CPU_wire_282_3,
CPU_wire_282_4,
CPU_wire_282_5,
CPU_wire_294_0,
CPU_wire_294_1,
CPU_wire_294_2,
CPU_wire_294_3,
CPU_wire_294_4,
CPU_wire_294_5,
CPU_wire_306_0,
CPU_wire_306_1,
CPU_wire_306_2,
CPU_wire_306_3,
CPU_wire_306_4,
CPU_wire_306_5,
CPU_wire_318_0,
CPU_wire_318_1,
CPU_wire_318_2,
CPU_wire_318_3,
CPU_wire_318_4,
CPU_wire_318_5,
CPU_wire_330_0,
CPU_wire_330_1,
CPU_wire_330_2,
CPU_wire_330_3,
CPU_wire_126_0,
CPU_wire_126_1,
CPU_wire_142_0,
CPU_wire_142_1,
CPU_wire_158_0,
CPU_wire_158_1,
CPU_wire_174_0,
CPU_wire_174_1,
CPU_wire_190_0,
CPU_wire_190_1,
CPU_wire_206_0,
CPU_wire_206_1,
CPU_wire_222_0,
CPU_wire_222_1,
CPU_wire_238_0,
CPU_wire_238_1,
CPU_wire_116_0,
CPU_wire_116_1,
CPU_wire_132_0,
CPU_wire_132_1,
CPU_wire_148_0,
CPU_wire_148_1,
CPU_wire_164_0,
CPU_wire_164_1,
CPU_wire_180_0,
CPU_wire_180_1,
CPU_wire_196_0,
CPU_wire_196_1,
CPU_wire_212_0,
CPU_wire_212_1,
CPU_wire_228_0,
CPU_wire_228_1,
CPU_wire_123_0,
CPU_wire_123_1,
CPU_wire_139_0,
CPU_wire_139_1,
CPU_wire_155_0,
CPU_wire_155_1,
CPU_wire_171_0,
CPU_wire_171_1,
CPU_wire_187_0,
CPU_wire_187_1,
CPU_wire_203_0,
CPU_wire_203_1,
CPU_wire_219_0,
CPU_wire_219_1,
CPU_wire_235_0,
CPU_wire_235_1,
CPU_wire_112_0,
CPU_wire_112_1,
CPU_wire_128_0,
CPU_wire_128_1,
CPU_wire_144_0,
CPU_wire_144_1,
CPU_wire_160_0,
CPU_wire_160_1,
CPU_wire_176_0,
CPU_wire_176_1,
CPU_wire_192_0,
CPU_wire_192_1,
CPU_wire_208_0,
CPU_wire_208_1,
CPU_wire_224_0,
CPU_wire_224_1,
CPU_wire_446_0,
CPU_wire_446_1,
CPU_wire_446_2,
CPU_wire_447_0,
CPU_wire_447_1,
CPU_wire_447_2,
CPU_wire_449_0,
CPU_wire_449_1,
CPU_wire_449_2,
CPU_wire_451_0,
CPU_wire_451_1,
CPU_wire_451_2,
CPU_wire_453_0,
CPU_wire_453_1,
CPU_wire_453_2,
CPU_wire_455_0,
CPU_wire_455_1,
CPU_wire_455_2,
CPU_wire_457_0,
CPU_wire_457_1,
CPU_wire_457_2,
CPU_wire_450_0,
CPU_wire_450_1,
CPU_wire_448_0,
CPU_wire_448_1,
CPU_wire_452_0,
CPU_wire_452_1,
CPU_wire_454_0,
CPU_wire_454_1,
CPU_wire_456_0,
CPU_wire_456_1,
CPU_wire_10_0,
CPU_wire_10_1,
CPU_wire_10_2,
CPU_wire_10_3,
CPU_wire_10_4,
CPU_wire_10_5,
CPU_wire_10_6,
CPU_wire_10_7,
CPU_wire_12_0,
CPU_wire_12_1,
CPU_wire_12_2,
CPU_wire_12_3,
CPU_wire_12_4,
CPU_wire_14_0,
CPU_wire_14_1,
CPU_wire_14_2,
CPU_wire_14_3,
CPU_wire_14_4,
CPU_wire_16_0,
CPU_wire_16_1,
CPU_wire_16_2,
CPU_wire_16_3,
CPU_wire_16_4,
CPU_wire_18_0,
CPU_wire_18_1,
CPU_wire_18_2,
CPU_wire_18_3,
CPU_wire_18_4,
CPU_wire_20_0,
CPU_wire_20_1,
CPU_wire_20_2,
CPU_wire_20_3,
CPU_wire_20_4,
CPU_wire_22_0,
CPU_wire_22_1,
CPU_wire_22_2,
CPU_wire_22_3,
CPU_wire_22_4,
CPU_wire_24_0,
CPU_wire_24_1,
CPU_wire_24_2,
CPU_wire_567_0,
CPU_wire_567_1,
CPU_wire_567_2,
CPU_wire_564_0,
CPU_wire_564_1,
CPU_wire_564_2,
CPU_wire_561_0,
CPU_wire_561_1,
CPU_wire_561_2,
CPU_wire_558_0,
CPU_wire_558_1,
CPU_wire_558_2,
CPU_wire_555_0,
CPU_wire_555_1,
CPU_wire_555_2,
CPU_wire_552_0,
CPU_wire_552_1,
CPU_wire_552_2,
CPU_wire_545_0,
CPU_wire_545_1,
CPU_wire_545_2,
CPU_wire_542_0,
CPU_wire_542_1,
CPU_wire_542_2,
CPU_wire_539_0,
CPU_wire_539_1,
CPU_wire_539_2,
CPU_wire_536_0,
CPU_wire_536_1,
CPU_wire_536_2,
CPU_wire_533_0,
CPU_wire_533_1,
CPU_wire_533_2,
CPU_wire_530_0,
CPU_wire_530_1,
CPU_wire_530_2,
CPU_wire_58_0,
CPU_wire_58_1,
CPU_wire_61_0,
CPU_wire_61_1,
CPU_wire_63_0,
CPU_wire_63_1,
CPU_wire_65_0,
CPU_wire_65_1,
CPU_wire_67_0,
CPU_wire_67_1,
CPU_wire_69_0,
CPU_wire_69_1,
CPU_wire_71_0,
CPU_wire_71_1,
CPU_wire_73_0,
CPU_wire_73_1,
CPU_wire_619_0,
CPU_wire_619_1,
CPU_wire_622_0,
CPU_wire_622_1,
CPU_wire_625_0,
CPU_wire_625_1,
CPU_wire_628_0,
CPU_wire_628_1,
CPU_wire_631_0,
CPU_wire_631_1,
CPU_wire_634_0,
CPU_wire_634_1,
CPU_wire_637_0,
CPU_wire_637_1,
CPU_wire_640_0,
CPU_wire_640_1,
CPU_wire_642_0,
CPU_wire_642_1,
CPU_wire_642_2,
CPU_wire_642_3,
CPU_wire_642_4,
CPU_wire_642_5,
CPU_wire_642_6,
CPU_wire_642_7,
CPU_wire_642_8,
CPU_wire_642_9,
CPU_wire_642_10,
CPU_wire_642_11,
CPU_wire_642_12,
CPU_wire_642_13,
CPU_wire_642_14,
CPU_wire_642_15,
CPU_wire_642_16,
CPU_wire_642_17,
CPU_wire_642_18,
CPU_wire_642_19,
CPU_wire_642_20,
CPU_wire_642_21,
CPU_wire_642_22,
CPU_wire_642_23,
CPU_wire_642_24,
CPU_wire_642_25,
CPU_wire_642_26,
CPU_wire_642_27,
CPU_wire_642_28,
CPU_wire_642_29,
CPU_wire_642_30,
CPU_wire_642_31,
CPU_wire_685_0,
CPU_wire_685_1,
CPU_wire_685_2,
CPU_wire_685_3,
CPU_wire_685_4,
CPU_wire_685_5,
CPU_wire_685_6,
CPU_wire_685_7,
CPU_wire_685_8,
CPU_wire_685_9,
CPU_wire_685_10,
CPU_wire_685_11,
CPU_wire_685_12,
CPU_wire_685_13,
CPU_wire_685_14,
CPU_wire_685_15,
CPU_wire_737_0,
CPU_wire_737_1,
CPU_wire_737_2,
CPU_wire_735_0,
CPU_wire_735_1,
CPU_wire_735_2,
CPU_wire_733_0,
CPU_wire_733_1,
CPU_wire_733_2,
CPU_wire_731_0,
CPU_wire_731_1,
CPU_wire_729_0,
CPU_wire_729_1,
CPU_wire_727_0,
CPU_wire_727_1,
CPU_wire_110_0,
CPU_wire_110_1,
CPU_wire_110_2,
CPU_wire_110_3,
CPU_wire_110_4,
CPU_wire_110_5,
CPU_wire_110_6,
CPU_wire_110_7,
CPU_wire_110_8,
CPU_wire_110_9,
CPU_wire_110_10,
CPU_wire_110_11,
CPU_wire_110_12,
CPU_wire_110_13,
CPU_wire_110_14,
CPU_wire_110_15,
CPU_wire_110_16,
CPU_wire_110_17,
CPU_wire_110_18,
CPU_wire_110_19,
clk_net_0,
reset_net_0,
store_net_0;
/* PPI0, PPI1, PPI2, PPI3, PPI4,PPI5, PPI6, PPI7, PPI8, PPI9,PPI10, PPI11, PPI12, PPI13, PPI14,PPI15, PPI16, PPI17, PPI18, PPI19,
PPI20, PPI21, PPI22, PPI23, PPI24,PPI25, PPI26, PPI27, PPI28, PPI29,PPI30, PPI31, PPI32, PPI33, PPI34,PPI35, PPI36, PPI37, PPI38, PPI39,
PPI40, PPI41, PPI42, PPI43, PPI44,PPI45, PPI46, PPI47, PPI48, PPI49,PPI50, PPI51, PPI52, PPI53, PPI54,PPI55,
PPO0, PPO1, PPO2, PPO3, PPO4,PPO5, PPO6, PPO7, PPO8, PPO9,PPO10, PPO11, PPO12, PPO13, PPO14,PPO15, PPO16, PPO17, PPO18, PPO19,
PPO20, PPO21, PPO22, PPO23, PPO24,PPO25, PPO26, PPO27, PPO28, PPO29,PPO30, PPO31, PPO32, PPO33, PPO34,PPO35, PPO36, PPO37, PPO38, PPO39,
PPO40, PPO41, PPO42, PPO43, PPO44,PPO45, PPO46, PPO47, PPO48, PPO49,PPO50, PPO51, PPO52, PPO53, PPO54,PPO55; */

pin #(8) pin_0 ({ inst[0], inst[1], inst[2], inst[3], inst[4], inst[5], inst[6], inst[7]}, {inst_0, inst_1, inst_2, inst_3, inst_4, inst_5, inst_6, inst_7});
//PPI

/* pin #(56) pin_1 ({CPU_wire_83,CPU_wire_84,CPU_wire_85,CPU_wire_87,CPU_wire_89,CPU_wire_90,CPU_wire_91,CPU_wire_93,
CPU_wire_337,CPU_wire_338,CPU_wire_339,CPU_wire_340,CPU_wire_341,CPU_wire_342,CPU_wire_343,CPU_wire_344,CPU_wire_346,CPU_wire_347,CPU_wire_348,CPU_wire_349,
CPU_wire_350,CPU_wire_351,CPU_wire_352,CPU_wire_353,CPU_wire_355,CPU_wire_356,CPU_wire_357,CPU_wire_358,CPU_wire_359,CPU_wire_360,CPU_wire_361,CPU_wire_362,
CPU_wire_364,CPU_wire_365,CPU_wire_366,CPU_wire_367,CPU_wire_368,CPU_wire_369,CPU_wire_370,CPU_wire_371,CPU_wire_501,CPU_wire_503,CPU_wire_505,CPU_wire_507,
CPU_wire_509,CPU_wire_511,CPU_wire_513,CPU_wire_515,CPU_wire_619,CPU_wire_622,CPU_wire_625,CPU_wire_628,CPU_wire_631,CPU_wire_634,CPU_wire_637,CPU_wire_640},
{PPI0, PPI1, PPI2, PPI3, PPI4,PPI5, PPI6, PPI7, PPI8, PPI9,PPI10, PPI11, PPI12, PPI13, PPI14,PPI15, PPI16, PPI17, PPI18, PPI19,
PPI20, PPI21, PPI22, PPI23, PPI24,PPI25, PPI26, PPI27, PPI28, PPI29,PPI30, PPI31, PPI32, PPI33, PPI34,PPI35, PPI36, PPI37, PPI38, PPI39,
PPI40, PPI41, PPI42, PPI43, PPI44,PPI45, PPI46, PPI47, PPI48, PPI49,PPI50, PPI51, PPI52, PPI53, PPI54,PPI55}); */


pout #(17) pout_0 ({address_0, address_1, address_2, address_3, address_4, address_5, address_6, address_7, out_data_0, out_data_1, out_data_2, out_data_3, out_data_4, out_data_5, out_data_6, out_data_7, store_net_0}, {address[0], address[1], address[2], address[3], address[4], address[5], address[6], address[7], out_data[0], out_data[1], out_data[2], out_data[3], out_data[4], out_data[5], out_data[6], out_data[7], store});

//PPO
/* pout #(56) pout_1 ({PPO0, PPO1, PPO2, PPO3, PPO4,PPO5, PPO6, PPO7, PPO8, PPO9,PPO10, PPO11, PPO12, PPO13, PPO14,PPO15, PPO16, PPO17, PPO18, PPO19,
PPO20, PPO21, PPO22, PPO23, PPO24,PPO25, PPO26, PPO27, PPO28, PPO29,PPO30, PPO31, PPO32, PPO33, PPO34,PPO35, PPO36, PPO37, PPO38, PPO39,
PPO40, PPO41, PPO42, PPO43, PPO44,PPO45, PPO46, PPO47, PPO48, PPO49,PPO50, PPO51, PPO52, PPO53, PPO54,PPO55},
{CPU_wire_75_outG,CPU_wire_78_outG,CPU_wire_86_outG,CPU_wire_88_outG,CPU_wire_2_outG,CPU_wire_4_outG,CPU_wire_92_outG,CPU_wire_7_outG,
CPU_wire_126_outG,CPU_wire_142_outG,CPU_wire_158_outG,CPU_wire_174_outG,CPU_wire_190_outG,CPU_wire_206_outG,CPU_wire_222_outG,CPU_wire_238_outG,CPU_wire_116_outG,
CPU_wire_132_outG,CPU_wire_148_outG,CPU_wire_164_outG,CPU_wire_180_outG,CPU_wire_196_outG, CPU_wire_212_outG,CPU_wire_228_outG,CPU_wire_123_outG,CPU_wire_139_outG,
CPU_wire_155_outG,CPU_wire_171_outG,CPU_wire_187_outG,CPU_wire_203_outG,CPU_wire_219_outG,CPU_wire_235_outG,CPU_wire_112_outG, CPU_wire_128_outG,CPU_wire_144_outG,
CPU_wire_160_outG,CPU_wire_176_outG,CPU_wire_192_outG,CPU_wire_208_outG,CPU_wire_224_outG,CPU_wire_10_outG,CPU_wire_12_outG,CPU_wire_14_outG,CPU_wire_16_outG,CPU_wire_18_outG,
CPU_wire_20_outG,CPU_wire_22_outG,CPU_wire_24_outG,CPU_wire_58_outG,CPU_wire_61_outG,CPU_wire_63_outG,CPU_wire_65_outG,CPU_wire_67_outG,
CPU_wire_69_outG,CPU_wire_71_outG,CPU_wire_73_outG}); */

fanout_n #(32, 0, 0) FANOUT_1 (CPU_wire_6, {CPU_wire_6_0, CPU_wire_6_1, CPU_wire_6_2, CPU_wire_6_3, CPU_wire_6_4, CPU_wire_6_5, CPU_wire_6_6, CPU_wire_6_7, CPU_wire_6_8, CPU_wire_6_9, CPU_wire_6_10, CPU_wire_6_11, CPU_wire_6_12, CPU_wire_6_13, CPU_wire_6_14, CPU_wire_6_15, CPU_wire_6_16, CPU_wire_6_17, CPU_wire_6_18, CPU_wire_6_19, CPU_wire_6_20, CPU_wire_6_21, CPU_wire_6_22, CPU_wire_6_23, CPU_wire_6_24, CPU_wire_6_25, CPU_wire_6_26, CPU_wire_6_27, CPU_wire_6_28, CPU_wire_6_29, CPU_wire_6_30, CPU_wire_6_31});
fanout_n #(36, 0, 0) FANOUT_2 (CPU_wire_8, {CPU_wire_8_0, CPU_wire_8_1, CPU_wire_8_2, CPU_wire_8_3, CPU_wire_8_4, CPU_wire_8_5, CPU_wire_8_6, CPU_wire_8_7, CPU_wire_8_8, CPU_wire_8_9, CPU_wire_8_10, CPU_wire_8_11, CPU_wire_8_12, CPU_wire_8_13, CPU_wire_8_14, CPU_wire_8_15, CPU_wire_8_16, CPU_wire_8_17, CPU_wire_8_18, CPU_wire_8_19, CPU_wire_8_20, CPU_wire_8_21, CPU_wire_8_22, CPU_wire_8_23, CPU_wire_8_24, CPU_wire_8_25, CPU_wire_8_26, CPU_wire_8_27, CPU_wire_8_28, CPU_wire_8_29, CPU_wire_8_30, CPU_wire_8_31, CPU_wire_8_32, CPU_wire_8_33, CPU_wire_8_34, CPU_wire_8_35});
fanout_n #(2, 0, 0) FANOUT_3 (CPU_wire_49, {CPU_wire_49_0, CPU_wire_49_1});
fanout_n #(2, 0, 0) FANOUT_4 (CPU_wire_50, {CPU_wire_50_0, CPU_wire_50_1});
fanout_n #(2, 0, 0) FANOUT_5 (CPU_wire_51, {CPU_wire_51_0, CPU_wire_51_1});
fanout_n #(2, 0, 0) FANOUT_6 (CPU_wire_52, {CPU_wire_52_0, CPU_wire_52_1});
fanout_n #(2, 0, 0) FANOUT_7 (CPU_wire_53, {CPU_wire_53_0, CPU_wire_53_1});
fanout_n #(2, 0, 0) FANOUT_8 (CPU_wire_54, {CPU_wire_54_0, CPU_wire_54_1});
fanout_n #(2, 0, 0) FANOUT_9 (CPU_wire_55, {CPU_wire_55_0, CPU_wire_55_1});
fanout_n #(2, 0, 0) FANOUT_10 (CPU_wire_56, {CPU_wire_56_0, CPU_wire_56_1});
fanout_n #(4, 0, 0) FANOUT_11 (CPU_wire_62, {CPU_wire_62_0, CPU_wire_62_1, CPU_wire_62_2, CPU_wire_62_3});
fanout_n #(4, 0, 0) FANOUT_12 (CPU_wire_64, {CPU_wire_64_0, CPU_wire_64_1, CPU_wire_64_2, CPU_wire_64_3});
fanout_n #(4, 0, 0) FANOUT_13 (CPU_wire_66, {CPU_wire_66_0, CPU_wire_66_1, CPU_wire_66_2, CPU_wire_66_3});
fanout_n #(4, 0, 0) FANOUT_14 (CPU_wire_68, {CPU_wire_68_0, CPU_wire_68_1, CPU_wire_68_2, CPU_wire_68_3});
fanout_n #(4, 0, 0) FANOUT_15 (CPU_wire_70, {CPU_wire_70_0, CPU_wire_70_1, CPU_wire_70_2, CPU_wire_70_3});
fanout_n #(4, 0, 0) FANOUT_16 (CPU_wire_72, {CPU_wire_72_0, CPU_wire_72_1, CPU_wire_72_2, CPU_wire_72_3});
fanout_n #(4, 0, 0) FANOUT_17 (CPU_wire_80, {CPU_wire_80_0, CPU_wire_80_1, CPU_wire_80_2, CPU_wire_80_3});
fanout_n #(4, 0, 0) FANOUT_18 (CPU_wire_81, {CPU_wire_81_0, CPU_wire_81_1, CPU_wire_81_2, CPU_wire_81_3});
fanout_n #(19, 0, 0) FANOUT_19 (CPU_wire_75, {CPU_wire_75_0, CPU_wire_75_1, CPU_wire_75_2, CPU_wire_75_3, CPU_wire_75_4, CPU_wire_75_5, CPU_wire_75_6, CPU_wire_75_7, CPU_wire_75_8, CPU_wire_75_9, CPU_wire_75_10, CPU_wire_75_11, CPU_wire_75_12, CPU_wire_75_13, CPU_wire_75_14, CPU_wire_75_15, CPU_wire_75_16, CPU_wire_75_17, CPU_wire_75_18});
fanout_n #(36, 0, 0) FANOUT_20 (CPU_wire_78, {CPU_wire_78_0, CPU_wire_78_1, CPU_wire_78_2, CPU_wire_78_3, CPU_wire_78_4, CPU_wire_78_5, CPU_wire_78_6, CPU_wire_78_7, CPU_wire_78_8, CPU_wire_78_9, CPU_wire_78_10, CPU_wire_78_11, CPU_wire_78_12, CPU_wire_78_13, CPU_wire_78_14, CPU_wire_78_15, CPU_wire_78_16, CPU_wire_78_17, CPU_wire_78_18, CPU_wire_78_19, CPU_wire_78_20, CPU_wire_78_21, CPU_wire_78_22, CPU_wire_78_23, CPU_wire_78_24, CPU_wire_78_25, CPU_wire_78_26, CPU_wire_78_27, CPU_wire_78_28, CPU_wire_78_29, CPU_wire_78_30, CPU_wire_78_31, CPU_wire_78_32, CPU_wire_78_33, CPU_wire_78_34, CPU_wire_78_35});
fanout_n #(55, 0, 0) FANOUT_21 (CPU_wire_86, {CPU_wire_86_0, CPU_wire_86_1, CPU_wire_86_2, CPU_wire_86_3, CPU_wire_86_4, CPU_wire_86_5, CPU_wire_86_6, CPU_wire_86_7, CPU_wire_86_8, CPU_wire_86_9, CPU_wire_86_10, CPU_wire_86_11, CPU_wire_86_12, CPU_wire_86_13, CPU_wire_86_14, CPU_wire_86_15, CPU_wire_86_16, CPU_wire_86_17, CPU_wire_86_18, CPU_wire_86_19, CPU_wire_86_20, CPU_wire_86_21, CPU_wire_86_22, CPU_wire_86_23, CPU_wire_86_24, CPU_wire_86_25, CPU_wire_86_26, CPU_wire_86_27, CPU_wire_86_28, CPU_wire_86_29, CPU_wire_86_30, CPU_wire_86_31, CPU_wire_86_32, CPU_wire_86_33, CPU_wire_86_34, CPU_wire_86_35, CPU_wire_86_36, CPU_wire_86_37, CPU_wire_86_38, CPU_wire_86_39, CPU_wire_86_40, CPU_wire_86_41, CPU_wire_86_42, CPU_wire_86_43, CPU_wire_86_44, CPU_wire_86_45, CPU_wire_86_46, CPU_wire_86_47, CPU_wire_86_48, CPU_wire_86_49, CPU_wire_86_50, CPU_wire_86_51, CPU_wire_86_52, CPU_wire_86_53, CPU_wire_86_54});
fanout_n #(71, 0, 0) FANOUT_22 (CPU_wire_88, {CPU_wire_88_0, CPU_wire_88_1, CPU_wire_88_2, CPU_wire_88_3, CPU_wire_88_4, CPU_wire_88_5, CPU_wire_88_6, CPU_wire_88_7, CPU_wire_88_8, CPU_wire_88_9, CPU_wire_88_10, CPU_wire_88_11, CPU_wire_88_12, CPU_wire_88_13, CPU_wire_88_14, CPU_wire_88_15, CPU_wire_88_16, CPU_wire_88_17, CPU_wire_88_18, CPU_wire_88_19, CPU_wire_88_20, CPU_wire_88_21, CPU_wire_88_22, CPU_wire_88_23, CPU_wire_88_24, CPU_wire_88_25, CPU_wire_88_26, CPU_wire_88_27, CPU_wire_88_28, CPU_wire_88_29, CPU_wire_88_30, CPU_wire_88_31, CPU_wire_88_32, CPU_wire_88_33, CPU_wire_88_34, CPU_wire_88_35, CPU_wire_88_36, CPU_wire_88_37, CPU_wire_88_38, CPU_wire_88_39, CPU_wire_88_40, CPU_wire_88_41, CPU_wire_88_42, CPU_wire_88_43, CPU_wire_88_44, CPU_wire_88_45, CPU_wire_88_46, CPU_wire_88_47, CPU_wire_88_48, CPU_wire_88_49, CPU_wire_88_50, CPU_wire_88_51, CPU_wire_88_52, CPU_wire_88_53, CPU_wire_88_54, CPU_wire_88_55, CPU_wire_88_56, CPU_wire_88_57, CPU_wire_88_58, CPU_wire_88_59, CPU_wire_88_60, CPU_wire_88_61, CPU_wire_88_62, CPU_wire_88_63, CPU_wire_88_64, CPU_wire_88_65, CPU_wire_88_66, CPU_wire_88_67, CPU_wire_88_68, CPU_wire_88_69, CPU_wire_88_70});
fanout_n #(12, 0, 0) FANOUT_23 (CPU_wire_2, {CPU_wire_2_0, CPU_wire_2_1, CPU_wire_2_2, CPU_wire_2_3, CPU_wire_2_4, CPU_wire_2_5, CPU_wire_2_6, CPU_wire_2_7, CPU_wire_2_8, CPU_wire_2_9, CPU_wire_2_10, CPU_wire_2_11});
fanout_n #(13, 0, 0) FANOUT_24 (CPU_wire_4, {CPU_wire_4_0, CPU_wire_4_1, CPU_wire_4_2, CPU_wire_4_3, CPU_wire_4_4, CPU_wire_4_5, CPU_wire_4_6, CPU_wire_4_7, CPU_wire_4_8, CPU_wire_4_9, CPU_wire_4_10, CPU_wire_4_11, CPU_wire_4_12});
fanout_n #(18, 0, 0) FANOUT_25 (CPU_wire_7, {CPU_wire_7_0, CPU_wire_7_1, CPU_wire_7_2, CPU_wire_7_3, CPU_wire_7_4, CPU_wire_7_5, CPU_wire_7_6, CPU_wire_7_7, CPU_wire_7_8, CPU_wire_7_9, CPU_wire_7_10, CPU_wire_7_11, CPU_wire_7_12, CPU_wire_7_13, CPU_wire_7_14, CPU_wire_7_15, CPU_wire_7_16, CPU_wire_7_17});
fanout_n #(3, 0, 0) FANOUT_26 (CPU_wire_120, {CPU_wire_120_0, CPU_wire_120_1, CPU_wire_120_2});
fanout_n #(7, 0, 0) FANOUT_27 (CPU_wire_136, {CPU_wire_136_0, CPU_wire_136_1, CPU_wire_136_2, CPU_wire_136_3, CPU_wire_136_4, CPU_wire_136_5, CPU_wire_136_6});
fanout_n #(5, 0, 0) FANOUT_28 (CPU_wire_152, {CPU_wire_152_0, CPU_wire_152_1, CPU_wire_152_2, CPU_wire_152_3, CPU_wire_152_4});
fanout_n #(5, 0, 0) FANOUT_29 (CPU_wire_168, {CPU_wire_168_0, CPU_wire_168_1, CPU_wire_168_2, CPU_wire_168_3, CPU_wire_168_4});
fanout_n #(5, 0, 0) FANOUT_30 (CPU_wire_184, {CPU_wire_184_0, CPU_wire_184_1, CPU_wire_184_2, CPU_wire_184_3, CPU_wire_184_4});
fanout_n #(5, 0, 0) FANOUT_31 (CPU_wire_200, {CPU_wire_200_0, CPU_wire_200_1, CPU_wire_200_2, CPU_wire_200_3, CPU_wire_200_4});
fanout_n #(5, 0, 0) FANOUT_32 (CPU_wire_216, {CPU_wire_216_0, CPU_wire_216_1, CPU_wire_216_2, CPU_wire_216_3, CPU_wire_216_4});
fanout_n #(5, 0, 0) FANOUT_33 (CPU_wire_232, {CPU_wire_232_0, CPU_wire_232_1, CPU_wire_232_2, CPU_wire_232_3, CPU_wire_232_4});
fanout_n #(2, 0, 0) FANOUT_34 (CPU_wire_246, {CPU_wire_246_0, CPU_wire_246_1});
fanout_n #(6, 0, 0) FANOUT_35 (CPU_wire_258, {CPU_wire_258_0, CPU_wire_258_1, CPU_wire_258_2, CPU_wire_258_3, CPU_wire_258_4, CPU_wire_258_5});
fanout_n #(6, 0, 0) FANOUT_36 (CPU_wire_270, {CPU_wire_270_0, CPU_wire_270_1, CPU_wire_270_2, CPU_wire_270_3, CPU_wire_270_4, CPU_wire_270_5});
fanout_n #(6, 0, 0) FANOUT_37 (CPU_wire_282, {CPU_wire_282_0, CPU_wire_282_1, CPU_wire_282_2, CPU_wire_282_3, CPU_wire_282_4, CPU_wire_282_5});
fanout_n #(6, 0, 0) FANOUT_38 (CPU_wire_294, {CPU_wire_294_0, CPU_wire_294_1, CPU_wire_294_2, CPU_wire_294_3, CPU_wire_294_4, CPU_wire_294_5});
fanout_n #(6, 0, 0) FANOUT_39 (CPU_wire_306, {CPU_wire_306_0, CPU_wire_306_1, CPU_wire_306_2, CPU_wire_306_3, CPU_wire_306_4, CPU_wire_306_5});
fanout_n #(6, 0, 0) FANOUT_40 (CPU_wire_318, {CPU_wire_318_0, CPU_wire_318_1, CPU_wire_318_2, CPU_wire_318_3, CPU_wire_318_4, CPU_wire_318_5});
fanout_n #(4, 0, 0) FANOUT_41 (CPU_wire_330, {CPU_wire_330_0, CPU_wire_330_1, CPU_wire_330_2, CPU_wire_330_3});
fanout_n #(2, 0, 0) FANOUT_42 (CPU_wire_126, {CPU_wire_126_0, CPU_wire_126_1});
fanout_n #(2, 0, 0) FANOUT_43 (CPU_wire_142, {CPU_wire_142_0, CPU_wire_142_1});
fanout_n #(2, 0, 0) FANOUT_44 (CPU_wire_158, {CPU_wire_158_0, CPU_wire_158_1});
fanout_n #(2, 0, 0) FANOUT_45 (CPU_wire_174, {CPU_wire_174_0, CPU_wire_174_1});
fanout_n #(2, 0, 0) FANOUT_46 (CPU_wire_190, {CPU_wire_190_0, CPU_wire_190_1});
fanout_n #(2, 0, 0) FANOUT_47 (CPU_wire_206, {CPU_wire_206_0, CPU_wire_206_1});
fanout_n #(2, 0, 0) FANOUT_48 (CPU_wire_222, {CPU_wire_222_0, CPU_wire_222_1});
fanout_n #(2, 0, 0) FANOUT_49 (CPU_wire_238, {CPU_wire_238_0, CPU_wire_238_1});
fanout_n #(2, 0, 0) FANOUT_50 (CPU_wire_116, {CPU_wire_116_0, CPU_wire_116_1});
fanout_n #(2, 0, 0) FANOUT_51 (CPU_wire_132, {CPU_wire_132_0, CPU_wire_132_1});
fanout_n #(2, 0, 0) FANOUT_52 (CPU_wire_148, {CPU_wire_148_0, CPU_wire_148_1});
fanout_n #(2, 0, 0) FANOUT_53 (CPU_wire_164, {CPU_wire_164_0, CPU_wire_164_1});
fanout_n #(2, 0, 0) FANOUT_54 (CPU_wire_180, {CPU_wire_180_0, CPU_wire_180_1});
fanout_n #(2, 0, 0) FANOUT_55 (CPU_wire_196, {CPU_wire_196_0, CPU_wire_196_1});
fanout_n #(2, 0, 0) FANOUT_56 (CPU_wire_212, {CPU_wire_212_0, CPU_wire_212_1});
fanout_n #(2, 0, 0) FANOUT_57 (CPU_wire_228, {CPU_wire_228_0, CPU_wire_228_1});
fanout_n #(2, 0, 0) FANOUT_58 (CPU_wire_123, {CPU_wire_123_0, CPU_wire_123_1});
fanout_n #(2, 0, 0) FANOUT_59 (CPU_wire_139, {CPU_wire_139_0, CPU_wire_139_1});
fanout_n #(2, 0, 0) FANOUT_60 (CPU_wire_155, {CPU_wire_155_0, CPU_wire_155_1});
fanout_n #(2, 0, 0) FANOUT_61 (CPU_wire_171, {CPU_wire_171_0, CPU_wire_171_1});
fanout_n #(2, 0, 0) FANOUT_62 (CPU_wire_187, {CPU_wire_187_0, CPU_wire_187_1});
fanout_n #(2, 0, 0) FANOUT_63 (CPU_wire_203, {CPU_wire_203_0, CPU_wire_203_1});
fanout_n #(2, 0, 0) FANOUT_64 (CPU_wire_219, {CPU_wire_219_0, CPU_wire_219_1});
fanout_n #(2, 0, 0) FANOUT_65 (CPU_wire_235, {CPU_wire_235_0, CPU_wire_235_1});
fanout_n #(2, 0, 0) FANOUT_66 (CPU_wire_112, {CPU_wire_112_0, CPU_wire_112_1});
fanout_n #(2, 0, 0) FANOUT_67 (CPU_wire_128, {CPU_wire_128_0, CPU_wire_128_1});
fanout_n #(2, 0, 0) FANOUT_68 (CPU_wire_144, {CPU_wire_144_0, CPU_wire_144_1});
fanout_n #(2, 0, 0) FANOUT_69 (CPU_wire_160, {CPU_wire_160_0, CPU_wire_160_1});
fanout_n #(2, 0, 0) FANOUT_70 (CPU_wire_176, {CPU_wire_176_0, CPU_wire_176_1});
fanout_n #(2, 0, 0) FANOUT_71 (CPU_wire_192, {CPU_wire_192_0, CPU_wire_192_1});
fanout_n #(2, 0, 0) FANOUT_72 (CPU_wire_208, {CPU_wire_208_0, CPU_wire_208_1});
fanout_n #(2, 0, 0) FANOUT_73 (CPU_wire_224, {CPU_wire_224_0, CPU_wire_224_1});
fanout_n #(3, 0, 0) FANOUT_74 (CPU_wire_446, {CPU_wire_446_0, CPU_wire_446_1, CPU_wire_446_2});
fanout_n #(3, 0, 0) FANOUT_75 (CPU_wire_447, {CPU_wire_447_0, CPU_wire_447_1, CPU_wire_447_2});
fanout_n #(3, 0, 0) FANOUT_76 (CPU_wire_449, {CPU_wire_449_0, CPU_wire_449_1, CPU_wire_449_2});
fanout_n #(3, 0, 0) FANOUT_77 (CPU_wire_451, {CPU_wire_451_0, CPU_wire_451_1, CPU_wire_451_2});
fanout_n #(3, 0, 0) FANOUT_78 (CPU_wire_453, {CPU_wire_453_0, CPU_wire_453_1, CPU_wire_453_2});
fanout_n #(3, 0, 0) FANOUT_79 (CPU_wire_455, {CPU_wire_455_0, CPU_wire_455_1, CPU_wire_455_2});
fanout_n #(3, 0, 0) FANOUT_80 (CPU_wire_457, {CPU_wire_457_0, CPU_wire_457_1, CPU_wire_457_2});
fanout_n #(2, 0, 0) FANOUT_81 (CPU_wire_450, {CPU_wire_450_0, CPU_wire_450_1});
fanout_n #(2, 0, 0) FANOUT_82 (CPU_wire_448, {CPU_wire_448_0, CPU_wire_448_1});
fanout_n #(2, 0, 0) FANOUT_83 (CPU_wire_452, {CPU_wire_452_0, CPU_wire_452_1});
fanout_n #(2, 0, 0) FANOUT_84 (CPU_wire_454, {CPU_wire_454_0, CPU_wire_454_1});
fanout_n #(2, 0, 0) FANOUT_85 (CPU_wire_456, {CPU_wire_456_0, CPU_wire_456_1});
fanout_n #(8, 0, 0) FANOUT_86 (CPU_wire_10, {CPU_wire_10_0, CPU_wire_10_1, CPU_wire_10_2, CPU_wire_10_3, CPU_wire_10_4, CPU_wire_10_5, CPU_wire_10_6, CPU_wire_10_7});
fanout_n #(5, 0, 0) FANOUT_87 (CPU_wire_12, {CPU_wire_12_0, CPU_wire_12_1, CPU_wire_12_2, CPU_wire_12_3, CPU_wire_12_4});
fanout_n #(5, 0, 0) FANOUT_88 (CPU_wire_14, {CPU_wire_14_0, CPU_wire_14_1, CPU_wire_14_2, CPU_wire_14_3, CPU_wire_14_4});
fanout_n #(5, 0, 0) FANOUT_89 (CPU_wire_16, {CPU_wire_16_0, CPU_wire_16_1, CPU_wire_16_2, CPU_wire_16_3, CPU_wire_16_4});
fanout_n #(5, 0, 0) FANOUT_90 (CPU_wire_18, {CPU_wire_18_0, CPU_wire_18_1, CPU_wire_18_2, CPU_wire_18_3, CPU_wire_18_4});
fanout_n #(5, 0, 0) FANOUT_91 (CPU_wire_20, {CPU_wire_20_0, CPU_wire_20_1, CPU_wire_20_2, CPU_wire_20_3, CPU_wire_20_4});
fanout_n #(5, 0, 0) FANOUT_92 (CPU_wire_22, {CPU_wire_22_0, CPU_wire_22_1, CPU_wire_22_2, CPU_wire_22_3, CPU_wire_22_4});
fanout_n #(3, 0, 0) FANOUT_93 (CPU_wire_24, {CPU_wire_24_0, CPU_wire_24_1, CPU_wire_24_2});
fanout_n #(3, 0, 0) FANOUT_94 (CPU_wire_567, {CPU_wire_567_0, CPU_wire_567_1, CPU_wire_567_2});
fanout_n #(3, 0, 0) FANOUT_95 (CPU_wire_564, {CPU_wire_564_0, CPU_wire_564_1, CPU_wire_564_2});
fanout_n #(3, 0, 0) FANOUT_96 (CPU_wire_561, {CPU_wire_561_0, CPU_wire_561_1, CPU_wire_561_2});
fanout_n #(3, 0, 0) FANOUT_97 (CPU_wire_558, {CPU_wire_558_0, CPU_wire_558_1, CPU_wire_558_2});
fanout_n #(3, 0, 0) FANOUT_98 (CPU_wire_555, {CPU_wire_555_0, CPU_wire_555_1, CPU_wire_555_2});
fanout_n #(3, 0, 0) FANOUT_99 (CPU_wire_552, {CPU_wire_552_0, CPU_wire_552_1, CPU_wire_552_2});
fanout_n #(3, 0, 0) FANOUT_100 (CPU_wire_545, {CPU_wire_545_0, CPU_wire_545_1, CPU_wire_545_2});
fanout_n #(3, 0, 0) FANOUT_101 (CPU_wire_542, {CPU_wire_542_0, CPU_wire_542_1, CPU_wire_542_2});
fanout_n #(3, 0, 0) FANOUT_102 (CPU_wire_539, {CPU_wire_539_0, CPU_wire_539_1, CPU_wire_539_2});
fanout_n #(3, 0, 0) FANOUT_103 (CPU_wire_536, {CPU_wire_536_0, CPU_wire_536_1, CPU_wire_536_2});
fanout_n #(3, 0, 0) FANOUT_104 (CPU_wire_533, {CPU_wire_533_0, CPU_wire_533_1, CPU_wire_533_2});
fanout_n #(3, 0, 0) FANOUT_105 (CPU_wire_530, {CPU_wire_530_0, CPU_wire_530_1, CPU_wire_530_2});
fanout_n #(2, 0, 0) FANOUT_106 (CPU_wire_58, {CPU_wire_58_0, CPU_wire_58_1});
fanout_n #(2, 0, 0) FANOUT_107 (CPU_wire_61, {CPU_wire_61_0, CPU_wire_61_1});
fanout_n #(2, 0, 0) FANOUT_108 (CPU_wire_63, {CPU_wire_63_0, CPU_wire_63_1});
fanout_n #(2, 0, 0) FANOUT_109 (CPU_wire_65, {CPU_wire_65_0, CPU_wire_65_1});
fanout_n #(2, 0, 0) FANOUT_110 (CPU_wire_67, {CPU_wire_67_0, CPU_wire_67_1});
fanout_n #(2, 0, 0) FANOUT_111 (CPU_wire_69, {CPU_wire_69_0, CPU_wire_69_1});
fanout_n #(2, 0, 0) FANOUT_112 (CPU_wire_71, {CPU_wire_71_0, CPU_wire_71_1});
fanout_n #(2, 0, 0) FANOUT_113 (CPU_wire_73, {CPU_wire_73_0, CPU_wire_73_1});
fanout_n #(2, 0, 0) FANOUT_114 (CPU_wire_619, {CPU_wire_619_0, CPU_wire_619_1});
fanout_n #(2, 0, 0) FANOUT_115 (CPU_wire_622, {CPU_wire_622_0, CPU_wire_622_1});
fanout_n #(2, 0, 0) FANOUT_116 (CPU_wire_625, {CPU_wire_625_0, CPU_wire_625_1});
fanout_n #(2, 0, 0) FANOUT_117 (CPU_wire_628, {CPU_wire_628_0, CPU_wire_628_1});
fanout_n #(2, 0, 0) FANOUT_118 (CPU_wire_631, {CPU_wire_631_0, CPU_wire_631_1});
fanout_n #(2, 0, 0) FANOUT_119 (CPU_wire_634, {CPU_wire_634_0, CPU_wire_634_1});
fanout_n #(2, 0, 0) FANOUT_120 (CPU_wire_637, {CPU_wire_637_0, CPU_wire_637_1});
fanout_n #(2, 0, 0) FANOUT_121 (CPU_wire_640, {CPU_wire_640_0, CPU_wire_640_1});
fanout_n #(32, 0, 0) FANOUT_122 (CPU_wire_642, {CPU_wire_642_0, CPU_wire_642_1, CPU_wire_642_2, CPU_wire_642_3, CPU_wire_642_4, CPU_wire_642_5, CPU_wire_642_6, CPU_wire_642_7, CPU_wire_642_8, CPU_wire_642_9, CPU_wire_642_10, CPU_wire_642_11, CPU_wire_642_12, CPU_wire_642_13, CPU_wire_642_14, CPU_wire_642_15, CPU_wire_642_16, CPU_wire_642_17, CPU_wire_642_18, CPU_wire_642_19, CPU_wire_642_20, CPU_wire_642_21, CPU_wire_642_22, CPU_wire_642_23, CPU_wire_642_24, CPU_wire_642_25, CPU_wire_642_26, CPU_wire_642_27, CPU_wire_642_28, CPU_wire_642_29, CPU_wire_642_30, CPU_wire_642_31});
fanout_n #(16, 0, 0) FANOUT_123 (CPU_wire_685, {CPU_wire_685_0, CPU_wire_685_1, CPU_wire_685_2, CPU_wire_685_3, CPU_wire_685_4, CPU_wire_685_5, CPU_wire_685_6, CPU_wire_685_7, CPU_wire_685_8, CPU_wire_685_9, CPU_wire_685_10, CPU_wire_685_11, CPU_wire_685_12, CPU_wire_685_13, CPU_wire_685_14, CPU_wire_685_15});
fanout_n #(3, 0, 0) FANOUT_124 (CPU_wire_737, {CPU_wire_737_0, CPU_wire_737_1, CPU_wire_737_2});
fanout_n #(3, 0, 0) FANOUT_125 (CPU_wire_735, {CPU_wire_735_0, CPU_wire_735_1, CPU_wire_735_2});
fanout_n #(3, 0, 0) FANOUT_126 (CPU_wire_733, {CPU_wire_733_0, CPU_wire_733_1, CPU_wire_733_2});
fanout_n #(2, 0, 0) FANOUT_127 (CPU_wire_731, {CPU_wire_731_0, CPU_wire_731_1});
fanout_n #(2, 0, 0) FANOUT_128 (CPU_wire_729, {CPU_wire_729_0, CPU_wire_729_1});
fanout_n #(2, 0, 0) FANOUT_129 (CPU_wire_727, {CPU_wire_727_0, CPU_wire_727_1});
fanout_n #(20, 0, 0) FANOUT_130 (CPU_wire_110, {CPU_wire_110_0, CPU_wire_110_1, CPU_wire_110_2, CPU_wire_110_3, CPU_wire_110_4, CPU_wire_110_5, CPU_wire_110_6, CPU_wire_110_7, CPU_wire_110_8, CPU_wire_110_9, CPU_wire_110_10, CPU_wire_110_11, CPU_wire_110_12, CPU_wire_110_13, CPU_wire_110_14, CPU_wire_110_15, CPU_wire_110_16, CPU_wire_110_17, CPU_wire_110_18, CPU_wire_110_19});


notg #(0, 0) NOT_1 (CPU_wire_1, CPU_wire_2_0);
and_n #(2, 0, 0) AND_1 (CPU_wire_3, {CPU_wire_4_0, CPU_wire_1});
notg #(0, 0) NOT_2 (CPU_wire_5, CPU_wire_4_1);
notg #(0, 0) NOT_3 (CPU_wire_6, CPU_wire_7_0);
or_n #(2, 0, 0) OR_1 (CPU_wire_8, {CPU_wire_7_1, CPU_wire_5});
and_n #(2, 0, 0) AND_2 (CPU_wire_9, {CPU_wire_10_0, CPU_wire_7_2});
and_n #(2, 0, 0) AND_3 (CPU_wire_11, {CPU_wire_12_0, CPU_wire_7_3});
and_n #(2, 0, 0) AND_4 (CPU_wire_13, {CPU_wire_14_0, CPU_wire_7_4});
and_n #(2, 0, 0) AND_5 (CPU_wire_15, {CPU_wire_16_0, CPU_wire_7_5});
and_n #(2, 0, 0) AND_6 (CPU_wire_17, {CPU_wire_18_0, CPU_wire_7_6});
and_n #(2, 0, 0) AND_7 (CPU_wire_19, {CPU_wire_20_0, CPU_wire_7_7});
and_n #(2, 0, 0) AND_8 (CPU_wire_21, {CPU_wire_22_0, CPU_wire_7_8});
and_n #(2, 0, 0) AND_9 (CPU_wire_23, {CPU_wire_24_0, CPU_wire_7_9});
and_n #(2, 0, 0) AND_10 (CPU_wire_25, {CPU_wire_26, CPU_wire_27});
and_n #(2, 0, 0) AND_11 (CPU_wire_28, {CPU_wire_29, CPU_wire_30});
and_n #(2, 0, 0) AND_12 (CPU_wire_31, {CPU_wire_32, CPU_wire_33});
and_n #(2, 0, 0) AND_13 (CPU_wire_34, {CPU_wire_35, CPU_wire_36});
and_n #(2, 0, 0) AND_14 (CPU_wire_37, {CPU_wire_38, CPU_wire_39});
and_n #(2, 0, 0) AND_15 (CPU_wire_40, {CPU_wire_41, CPU_wire_42});
and_n #(2, 0, 0) AND_16 (CPU_wire_43, {CPU_wire_44, CPU_wire_45});
and_n #(2, 0, 0) AND_17 (CPU_wire_46, {CPU_wire_47, CPU_wire_48});
or_n #(2, 0, 0) OR_2 (CPU_wire_49, {CPU_wire_9, CPU_wire_25});
notg #(0, 0) NOT_4 (CPU_wire_27, CPU_wire_7_10);
or_n #(2, 0, 0) OR_3 (CPU_wire_50, {CPU_wire_11, CPU_wire_28});
notg #(0, 0) NOT_5 (CPU_wire_30, CPU_wire_7_11);
or_n #(2, 0, 0) OR_4 (CPU_wire_51, {CPU_wire_13, CPU_wire_31});
notg #(0, 0) NOT_6 (CPU_wire_33, CPU_wire_7_12);
or_n #(2, 0, 0) OR_5 (CPU_wire_52, {CPU_wire_15, CPU_wire_34});
notg #(0, 0) NOT_7 (CPU_wire_36, CPU_wire_7_13);
or_n #(2, 0, 0) OR_6 (CPU_wire_53, {CPU_wire_17, CPU_wire_37});
notg #(0, 0) NOT_8 (CPU_wire_39, CPU_wire_7_14);
or_n #(2, 0, 0) OR_7 (CPU_wire_54, {CPU_wire_19, CPU_wire_40});
notg #(0, 0) NOT_9 (CPU_wire_42, CPU_wire_7_15);
or_n #(2, 0, 0) OR_8 (CPU_wire_55, {CPU_wire_21, CPU_wire_43});
notg #(0, 0) NOT_10 (CPU_wire_45, CPU_wire_7_16);
or_n #(2, 0, 0) OR_9 (CPU_wire_56, {CPU_wire_23, CPU_wire_46});
notg #(0, 0) NOT_11 (CPU_wire_48, CPU_wire_7_17);
and_n #(2, 0, 0) AND_18 (CPU_wire_57, {CPU_wire_58_0, CPU_wire_59});
and_n #(2, 0, 0) AND_19 (CPU_wire_60, {CPU_wire_61_0, CPU_wire_59});
and_n #(2, 0, 0) AND_20 (CPU_wire_62, {CPU_wire_63_0, CPU_wire_59});
and_n #(2, 0, 0) AND_21 (CPU_wire_64, {CPU_wire_65_0, CPU_wire_59});
and_n #(2, 0, 0) AND_22 (CPU_wire_66, {CPU_wire_67_0, CPU_wire_59});
and_n #(2, 0, 0) AND_23 (CPU_wire_68, {CPU_wire_69_0, CPU_wire_59});
and_n #(2, 0, 0) AND_24 (CPU_wire_70, {CPU_wire_71_0, CPU_wire_59});
and_n #(2, 0, 0) AND_25 (CPU_wire_72, {CPU_wire_73_0, CPU_wire_59});
and_n #(2, 0, 0) AND_26 (CPU_wire_74, {CPU_wire_75_0, CPU_wire_76});
and_n #(2, 0, 0) AND_27 (CPU_wire_77, {CPU_wire_78_0, CPU_wire_79});
or_n #(2, 0, 0) OR_10 (CPU_wire_80, {CPU_wire_57, CPU_wire_74});
notg #(0, 0) NOT_12 (CPU_wire_76, CPU_wire_59);
or_n #(2, 0, 0) OR_11 (CPU_wire_81, {CPU_wire_60, CPU_wire_77});
notg #(0, 0) NOT_13 (CPU_wire_79, CPU_wire_59);
and_n #(2, 0, 0) AND_28 (CPU_wire_83, {CPU_wire_94, CPU_wire_95});
and_n #(2, 0, 0) AND_29 (CPU_wire_84, {CPU_wire_96, CPU_wire_97});
and_n #(2, 0, 0) AND_30 (CPU_wire_85, {CPU_wire_98, CPU_wire_99});
and_n #(2, 0, 0) AND_31 (CPU_wire_87, {CPU_wire_100, CPU_wire_101});
and_n #(2, 0, 0) AND_32 (CPU_wire_89, {CPU_wire_102, CPU_wire_103});
and_n #(2, 0, 0) AND_33 (CPU_wire_90, {CPU_wire_104, CPU_wire_105});
and_n #(2, 0, 0) AND_34 (CPU_wire_91, {CPU_wire_106, CPU_wire_107});
and_n #(2, 0, 0) AND_35 (CPU_wire_93, {CPU_wire_108, CPU_wire_109});
notg #(0, 0) NOT_14 (CPU_wire_95, CPU_wire_110_0);
notg #(0, 0) NOT_15 (CPU_wire_97, CPU_wire_110_1);
notg #(0, 0) NOT_16 (CPU_wire_99, CPU_wire_110_2);
notg #(0, 0) NOT_17 (CPU_wire_101, CPU_wire_110_3);
notg #(0, 0) NOT_18 (CPU_wire_103, CPU_wire_110_4);
notg #(0, 0) NOT_19 (CPU_wire_105, CPU_wire_110_5);
notg #(0, 0) NOT_20 (CPU_wire_107, CPU_wire_110_6);
notg #(0, 0) NOT_21 (CPU_wire_109, CPU_wire_110_7);
and_n #(2, 0, 0) AND_36 (CPU_wire_111, {CPU_wire_88_0, CPU_wire_112_0});
or_n #(2, 0, 0) OR_12 (CPU_wire_113, {CPU_wire_111, CPU_wire_114});
notg #(0, 0) NOT_22 (CPU_wire_115, CPU_wire_88_1);
and_n #(2, 0, 0) AND_37 (CPU_wire_114, {CPU_wire_115, CPU_wire_116_0});
and_n #(2, 0, 0) AND_38 (CPU_wire_117, {CPU_wire_118, CPU_wire_119});
or_n #(2, 0, 0) OR_13 (CPU_wire_120, {CPU_wire_117, CPU_wire_121});
and_n #(2, 0, 0) AND_39 (CPU_wire_122, {CPU_wire_88_2, CPU_wire_123_0});
or_n #(2, 0, 0) OR_14 (CPU_wire_119, {CPU_wire_122, CPU_wire_124});
notg #(0, 0) NOT_23 (CPU_wire_125, CPU_wire_88_3);
and_n #(2, 0, 0) AND_40 (CPU_wire_124, {CPU_wire_125, CPU_wire_126_0});
notg #(0, 0) NOT_24 (CPU_wire_118, CPU_wire_86_0);
and_n #(2, 0, 0) AND_41 (CPU_wire_121, {CPU_wire_113, CPU_wire_86_1});
and_n #(2, 0, 0) AND_42 (CPU_wire_127, {CPU_wire_88_4, CPU_wire_128_0});
or_n #(2, 0, 0) OR_15 (CPU_wire_129, {CPU_wire_127, CPU_wire_130});
notg #(0, 0) NOT_25 (CPU_wire_131, CPU_wire_88_5);
and_n #(2, 0, 0) AND_43 (CPU_wire_130, {CPU_wire_131, CPU_wire_132_0});
and_n #(2, 0, 0) AND_44 (CPU_wire_133, {CPU_wire_134, CPU_wire_135});
or_n #(2, 0, 0) OR_16 (CPU_wire_136, {CPU_wire_133, CPU_wire_137});
and_n #(2, 0, 0) AND_45 (CPU_wire_138, {CPU_wire_88_6, CPU_wire_139_0});
or_n #(2, 0, 0) OR_17 (CPU_wire_135, {CPU_wire_138, CPU_wire_140});
notg #(0, 0) NOT_26 (CPU_wire_141, CPU_wire_88_7);
and_n #(2, 0, 0) AND_46 (CPU_wire_140, {CPU_wire_141, CPU_wire_142_0});
notg #(0, 0) NOT_27 (CPU_wire_134, CPU_wire_86_2);
and_n #(2, 0, 0) AND_47 (CPU_wire_137, {CPU_wire_129, CPU_wire_86_3});
and_n #(2, 0, 0) AND_48 (CPU_wire_143, {CPU_wire_88_8, CPU_wire_144_0});
or_n #(2, 0, 0) OR_18 (CPU_wire_145, {CPU_wire_143, CPU_wire_146});
notg #(0, 0) NOT_28 (CPU_wire_147, CPU_wire_88_9);
and_n #(2, 0, 0) AND_49 (CPU_wire_146, {CPU_wire_147, CPU_wire_148_0});
and_n #(2, 0, 0) AND_50 (CPU_wire_149, {CPU_wire_150, CPU_wire_151});
or_n #(2, 0, 0) OR_19 (CPU_wire_152, {CPU_wire_149, CPU_wire_153});
and_n #(2, 0, 0) AND_51 (CPU_wire_154, {CPU_wire_88_10, CPU_wire_155_0});
or_n #(2, 0, 0) OR_20 (CPU_wire_151, {CPU_wire_154, CPU_wire_156});
notg #(0, 0) NOT_29 (CPU_wire_157, CPU_wire_88_11);
and_n #(2, 0, 0) AND_52 (CPU_wire_156, {CPU_wire_157, CPU_wire_158_0});
notg #(0, 0) NOT_30 (CPU_wire_150, CPU_wire_86_4);
and_n #(2, 0, 0) AND_53 (CPU_wire_153, {CPU_wire_145, CPU_wire_86_5});
and_n #(2, 0, 0) AND_54 (CPU_wire_159, {CPU_wire_88_12, CPU_wire_160_0});
or_n #(2, 0, 0) OR_21 (CPU_wire_161, {CPU_wire_159, CPU_wire_162});
notg #(0, 0) NOT_31 (CPU_wire_163, CPU_wire_88_13);
and_n #(2, 0, 0) AND_55 (CPU_wire_162, {CPU_wire_163, CPU_wire_164_0});
and_n #(2, 0, 0) AND_56 (CPU_wire_165, {CPU_wire_166, CPU_wire_167});
or_n #(2, 0, 0) OR_22 (CPU_wire_168, {CPU_wire_165, CPU_wire_169});
and_n #(2, 0, 0) AND_57 (CPU_wire_170, {CPU_wire_88_14, CPU_wire_171_0});
or_n #(2, 0, 0) OR_23 (CPU_wire_167, {CPU_wire_170, CPU_wire_172});
notg #(0, 0) NOT_32 (CPU_wire_173, CPU_wire_88_15);
and_n #(2, 0, 0) AND_58 (CPU_wire_172, {CPU_wire_173, CPU_wire_174_0});
notg #(0, 0) NOT_33 (CPU_wire_166, CPU_wire_86_6);
and_n #(2, 0, 0) AND_59 (CPU_wire_169, {CPU_wire_161, CPU_wire_86_7});
and_n #(2, 0, 0) AND_60 (CPU_wire_175, {CPU_wire_88_16, CPU_wire_176_0});
or_n #(2, 0, 0) OR_24 (CPU_wire_177, {CPU_wire_175, CPU_wire_178});
notg #(0, 0) NOT_34 (CPU_wire_179, CPU_wire_88_17);
and_n #(2, 0, 0) AND_61 (CPU_wire_178, {CPU_wire_179, CPU_wire_180_0});
and_n #(2, 0, 0) AND_62 (CPU_wire_181, {CPU_wire_182, CPU_wire_183});
or_n #(2, 0, 0) OR_25 (CPU_wire_184, {CPU_wire_181, CPU_wire_185});
and_n #(2, 0, 0) AND_63 (CPU_wire_186, {CPU_wire_88_18, CPU_wire_187_0});
or_n #(2, 0, 0) OR_26 (CPU_wire_183, {CPU_wire_186, CPU_wire_188});
notg #(0, 0) NOT_35 (CPU_wire_189, CPU_wire_88_19);
and_n #(2, 0, 0) AND_64 (CPU_wire_188, {CPU_wire_189, CPU_wire_190_0});
notg #(0, 0) NOT_36 (CPU_wire_182, CPU_wire_86_8);
and_n #(2, 0, 0) AND_65 (CPU_wire_185, {CPU_wire_177, CPU_wire_86_9});
and_n #(2, 0, 0) AND_66 (CPU_wire_191, {CPU_wire_88_20, CPU_wire_192_0});
or_n #(2, 0, 0) OR_27 (CPU_wire_193, {CPU_wire_191, CPU_wire_194});
notg #(0, 0) NOT_37 (CPU_wire_195, CPU_wire_88_21);
and_n #(2, 0, 0) AND_67 (CPU_wire_194, {CPU_wire_195, CPU_wire_196_0});
and_n #(2, 0, 0) AND_68 (CPU_wire_197, {CPU_wire_198, CPU_wire_199});
or_n #(2, 0, 0) OR_28 (CPU_wire_200, {CPU_wire_197, CPU_wire_201});
and_n #(2, 0, 0) AND_69 (CPU_wire_202, {CPU_wire_88_22, CPU_wire_203_0});
or_n #(2, 0, 0) OR_29 (CPU_wire_199, {CPU_wire_202, CPU_wire_204});
notg #(0, 0) NOT_38 (CPU_wire_205, CPU_wire_88_23);
and_n #(2, 0, 0) AND_70 (CPU_wire_204, {CPU_wire_205, CPU_wire_206_0});
notg #(0, 0) NOT_39 (CPU_wire_198, CPU_wire_86_10);
and_n #(2, 0, 0) AND_71 (CPU_wire_201, {CPU_wire_193, CPU_wire_86_11});
and_n #(2, 0, 0) AND_72 (CPU_wire_207, {CPU_wire_88_24, CPU_wire_208_0});
or_n #(2, 0, 0) OR_30 (CPU_wire_209, {CPU_wire_207, CPU_wire_210});
notg #(0, 0) NOT_40 (CPU_wire_211, CPU_wire_88_25);
and_n #(2, 0, 0) AND_73 (CPU_wire_210, {CPU_wire_211, CPU_wire_212_0});
and_n #(2, 0, 0) AND_74 (CPU_wire_213, {CPU_wire_214, CPU_wire_215});
or_n #(2, 0, 0) OR_31 (CPU_wire_216, {CPU_wire_213, CPU_wire_217});
and_n #(2, 0, 0) AND_75 (CPU_wire_218, {CPU_wire_88_26, CPU_wire_219_0});
or_n #(2, 0, 0) OR_32 (CPU_wire_215, {CPU_wire_218, CPU_wire_220});
notg #(0, 0) NOT_41 (CPU_wire_221, CPU_wire_88_27);
and_n #(2, 0, 0) AND_76 (CPU_wire_220, {CPU_wire_221, CPU_wire_222_0});
notg #(0, 0) NOT_42 (CPU_wire_214, CPU_wire_86_12);
and_n #(2, 0, 0) AND_77 (CPU_wire_217, {CPU_wire_209, CPU_wire_86_13});
and_n #(2, 0, 0) AND_78 (CPU_wire_223, {CPU_wire_88_28, CPU_wire_224_0});
or_n #(2, 0, 0) OR_33 (CPU_wire_225, {CPU_wire_223, CPU_wire_226});
notg #(0, 0) NOT_43 (CPU_wire_227, CPU_wire_88_29);
and_n #(2, 0, 0) AND_79 (CPU_wire_226, {CPU_wire_227, CPU_wire_228_0});
and_n #(2, 0, 0) AND_80 (CPU_wire_229, {CPU_wire_230, CPU_wire_231});
or_n #(2, 0, 0) OR_34 (CPU_wire_232, {CPU_wire_229, CPU_wire_233});
and_n #(2, 0, 0) AND_81 (CPU_wire_234, {CPU_wire_88_30, CPU_wire_235_0});
or_n #(2, 0, 0) OR_35 (CPU_wire_231, {CPU_wire_234, CPU_wire_236});
notg #(0, 0) NOT_44 (CPU_wire_237, CPU_wire_88_31);
and_n #(2, 0, 0) AND_82 (CPU_wire_236, {CPU_wire_237, CPU_wire_238_0});
notg #(0, 0) NOT_45 (CPU_wire_230, CPU_wire_86_14);
and_n #(2, 0, 0) AND_83 (CPU_wire_233, {CPU_wire_225, CPU_wire_86_15});
and_n #(2, 0, 0) AND_84 (CPU_wire_239, {CPU_wire_78_1, CPU_wire_112_1});
or_n #(2, 0, 0) OR_36 (CPU_wire_240, {CPU_wire_239, CPU_wire_241});
notg #(0, 0) NOT_46 (CPU_wire_242, CPU_wire_78_2);
and_n #(2, 0, 0) AND_85 (CPU_wire_241, {CPU_wire_242, CPU_wire_116_1});
and_n #(2, 0, 0) AND_86 (CPU_wire_243, {CPU_wire_244, CPU_wire_245});
or_n #(2, 0, 0) OR_37 (CPU_wire_246, {CPU_wire_243, CPU_wire_247});
and_n #(2, 0, 0) AND_87 (CPU_wire_248, {CPU_wire_78_3, CPU_wire_123_1});
or_n #(2, 0, 0) OR_38 (CPU_wire_245, {CPU_wire_248, CPU_wire_249});
notg #(0, 0) NOT_47 (CPU_wire_250, CPU_wire_78_4);
and_n #(2, 0, 0) AND_88 (CPU_wire_249, {CPU_wire_250, CPU_wire_126_1});
notg #(0, 0) NOT_48 (CPU_wire_244, CPU_wire_75_1);
and_n #(2, 0, 0) AND_89 (CPU_wire_247, {CPU_wire_240, CPU_wire_75_2});
and_n #(2, 0, 0) AND_90 (CPU_wire_251, {CPU_wire_78_5, CPU_wire_128_1});
or_n #(2, 0, 0) OR_39 (CPU_wire_252, {CPU_wire_251, CPU_wire_253});
notg #(0, 0) NOT_49 (CPU_wire_254, CPU_wire_78_6);
and_n #(2, 0, 0) AND_91 (CPU_wire_253, {CPU_wire_254, CPU_wire_132_1});
and_n #(2, 0, 0) AND_92 (CPU_wire_255, {CPU_wire_256, CPU_wire_257});
or_n #(2, 0, 0) OR_40 (CPU_wire_258, {CPU_wire_255, CPU_wire_259});
and_n #(2, 0, 0) AND_93 (CPU_wire_260, {CPU_wire_78_7, CPU_wire_139_1});
or_n #(2, 0, 0) OR_41 (CPU_wire_257, {CPU_wire_260, CPU_wire_261});
notg #(0, 0) NOT_50 (CPU_wire_262, CPU_wire_78_8);
and_n #(2, 0, 0) AND_94 (CPU_wire_261, {CPU_wire_262, CPU_wire_142_1});
notg #(0, 0) NOT_51 (CPU_wire_256, CPU_wire_75_3);
and_n #(2, 0, 0) AND_95 (CPU_wire_259, {CPU_wire_252, CPU_wire_75_4});
and_n #(2, 0, 0) AND_96 (CPU_wire_263, {CPU_wire_78_9, CPU_wire_144_1});
or_n #(2, 0, 0) OR_42 (CPU_wire_264, {CPU_wire_263, CPU_wire_265});
notg #(0, 0) NOT_52 (CPU_wire_266, CPU_wire_78_10);
and_n #(2, 0, 0) AND_97 (CPU_wire_265, {CPU_wire_266, CPU_wire_148_1});
and_n #(2, 0, 0) AND_98 (CPU_wire_267, {CPU_wire_268, CPU_wire_269});
or_n #(2, 0, 0) OR_43 (CPU_wire_270, {CPU_wire_267, CPU_wire_271});
and_n #(2, 0, 0) AND_99 (CPU_wire_272, {CPU_wire_78_11, CPU_wire_155_1});
or_n #(2, 0, 0) OR_44 (CPU_wire_269, {CPU_wire_272, CPU_wire_273});
notg #(0, 0) NOT_53 (CPU_wire_274, CPU_wire_78_12);
and_n #(2, 0, 0) AND_100 (CPU_wire_273, {CPU_wire_274, CPU_wire_158_1});
notg #(0, 0) NOT_54 (CPU_wire_268, CPU_wire_75_5);
and_n #(2, 0, 0) AND_101 (CPU_wire_271, {CPU_wire_264, CPU_wire_75_6});
and_n #(2, 0, 0) AND_102 (CPU_wire_275, {CPU_wire_78_13, CPU_wire_160_1});
or_n #(2, 0, 0) OR_45 (CPU_wire_276, {CPU_wire_275, CPU_wire_277});
notg #(0, 0) NOT_55 (CPU_wire_278, CPU_wire_78_14);
and_n #(2, 0, 0) AND_103 (CPU_wire_277, {CPU_wire_278, CPU_wire_164_1});
and_n #(2, 0, 0) AND_104 (CPU_wire_279, {CPU_wire_280, CPU_wire_281});
or_n #(2, 0, 0) OR_46 (CPU_wire_282, {CPU_wire_279, CPU_wire_283});
and_n #(2, 0, 0) AND_105 (CPU_wire_284, {CPU_wire_78_15, CPU_wire_171_1});
or_n #(2, 0, 0) OR_47 (CPU_wire_281, {CPU_wire_284, CPU_wire_285});
notg #(0, 0) NOT_56 (CPU_wire_286, CPU_wire_78_16);
and_n #(2, 0, 0) AND_106 (CPU_wire_285, {CPU_wire_286, CPU_wire_174_1});
notg #(0, 0) NOT_57 (CPU_wire_280, CPU_wire_75_7);
and_n #(2, 0, 0) AND_107 (CPU_wire_283, {CPU_wire_276, CPU_wire_75_8});
and_n #(2, 0, 0) AND_108 (CPU_wire_287, {CPU_wire_78_17, CPU_wire_176_1});
or_n #(2, 0, 0) OR_48 (CPU_wire_288, {CPU_wire_287, CPU_wire_289});
notg #(0, 0) NOT_58 (CPU_wire_290, CPU_wire_78_18);
and_n #(2, 0, 0) AND_109 (CPU_wire_289, {CPU_wire_290, CPU_wire_180_1});
and_n #(2, 0, 0) AND_110 (CPU_wire_291, {CPU_wire_292, CPU_wire_293});
or_n #(2, 0, 0) OR_49 (CPU_wire_294, {CPU_wire_291, CPU_wire_295});
and_n #(2, 0, 0) AND_111 (CPU_wire_296, {CPU_wire_78_19, CPU_wire_187_1});
or_n #(2, 0, 0) OR_50 (CPU_wire_293, {CPU_wire_296, CPU_wire_297});
notg #(0, 0) NOT_59 (CPU_wire_298, CPU_wire_78_20);
and_n #(2, 0, 0) AND_112 (CPU_wire_297, {CPU_wire_298, CPU_wire_190_1});
notg #(0, 0) NOT_60 (CPU_wire_292, CPU_wire_75_9);
and_n #(2, 0, 0) AND_113 (CPU_wire_295, {CPU_wire_288, CPU_wire_75_10});
and_n #(2, 0, 0) AND_114 (CPU_wire_299, {CPU_wire_78_21, CPU_wire_192_1});
or_n #(2, 0, 0) OR_51 (CPU_wire_300, {CPU_wire_299, CPU_wire_301});
notg #(0, 0) NOT_61 (CPU_wire_302, CPU_wire_78_22);
and_n #(2, 0, 0) AND_115 (CPU_wire_301, {CPU_wire_302, CPU_wire_196_1});
and_n #(2, 0, 0) AND_116 (CPU_wire_303, {CPU_wire_304, CPU_wire_305});
or_n #(2, 0, 0) OR_52 (CPU_wire_306, {CPU_wire_303, CPU_wire_307});
and_n #(2, 0, 0) AND_117 (CPU_wire_308, {CPU_wire_78_23, CPU_wire_203_1});
or_n #(2, 0, 0) OR_53 (CPU_wire_305, {CPU_wire_308, CPU_wire_309});
notg #(0, 0) NOT_62 (CPU_wire_310, CPU_wire_78_24);
and_n #(2, 0, 0) AND_118 (CPU_wire_309, {CPU_wire_310, CPU_wire_206_1});
notg #(0, 0) NOT_63 (CPU_wire_304, CPU_wire_75_11);
and_n #(2, 0, 0) AND_119 (CPU_wire_307, {CPU_wire_300, CPU_wire_75_12});
and_n #(2, 0, 0) AND_120 (CPU_wire_311, {CPU_wire_78_25, CPU_wire_208_1});
or_n #(2, 0, 0) OR_54 (CPU_wire_312, {CPU_wire_311, CPU_wire_313});
notg #(0, 0) NOT_64 (CPU_wire_314, CPU_wire_78_26);
and_n #(2, 0, 0) AND_121 (CPU_wire_313, {CPU_wire_314, CPU_wire_212_1});
and_n #(2, 0, 0) AND_122 (CPU_wire_315, {CPU_wire_316, CPU_wire_317});
or_n #(2, 0, 0) OR_55 (CPU_wire_318, {CPU_wire_315, CPU_wire_319});
and_n #(2, 0, 0) AND_123 (CPU_wire_320, {CPU_wire_78_27, CPU_wire_219_1});
or_n #(2, 0, 0) OR_56 (CPU_wire_317, {CPU_wire_320, CPU_wire_321});
notg #(0, 0) NOT_65 (CPU_wire_322, CPU_wire_78_28);
and_n #(2, 0, 0) AND_124 (CPU_wire_321, {CPU_wire_322, CPU_wire_222_1});
notg #(0, 0) NOT_66 (CPU_wire_316, CPU_wire_75_13);
and_n #(2, 0, 0) AND_125 (CPU_wire_319, {CPU_wire_312, CPU_wire_75_14});
and_n #(2, 0, 0) AND_126 (CPU_wire_323, {CPU_wire_78_29, CPU_wire_224_1});
or_n #(2, 0, 0) OR_57 (CPU_wire_324, {CPU_wire_323, CPU_wire_325});
notg #(0, 0) NOT_67 (CPU_wire_326, CPU_wire_78_30);
and_n #(2, 0, 0) AND_127 (CPU_wire_325, {CPU_wire_326, CPU_wire_228_1});
and_n #(2, 0, 0) AND_128 (CPU_wire_327, {CPU_wire_328, CPU_wire_329});
or_n #(2, 0, 0) OR_58 (CPU_wire_330, {CPU_wire_327, CPU_wire_331});
and_n #(2, 0, 0) AND_129 (CPU_wire_332, {CPU_wire_78_31, CPU_wire_235_1});
or_n #(2, 0, 0) OR_59 (CPU_wire_329, {CPU_wire_332, CPU_wire_333});
notg #(0, 0) NOT_68 (CPU_wire_334, CPU_wire_78_32);
and_n #(2, 0, 0) AND_130 (CPU_wire_333, {CPU_wire_334, CPU_wire_238_1});
notg #(0, 0) NOT_69 (CPU_wire_328, CPU_wire_75_15);
and_n #(2, 0, 0) AND_131 (CPU_wire_331, {CPU_wire_324, CPU_wire_75_16});
bufg #(0, 0) BUF_1 (CPU_wire_335, 1'b0);
and_n #(2, 0, 0) AND_132 (CPU_wire_372, {CPU_wire_86_16, CPU_wire_373});
and_n #(2, 0, 0) AND_133 (CPU_wire_374, {CPU_wire_86_17, CPU_wire_375});
and_n #(2, 0, 0) AND_134 (CPU_wire_376, {CPU_wire_86_18, CPU_wire_377});
and_n #(2, 0, 0) AND_135 (CPU_wire_378, {CPU_wire_86_19, CPU_wire_379});
and_n #(2, 0, 0) AND_136 (CPU_wire_380, {CPU_wire_86_20, CPU_wire_381});
and_n #(2, 0, 0) AND_137 (CPU_wire_382, {CPU_wire_86_21, CPU_wire_383});
and_n #(2, 0, 0) AND_138 (CPU_wire_384, {CPU_wire_86_22, CPU_wire_385});
and_n #(2, 0, 0) AND_139 (CPU_wire_386, {CPU_wire_86_23, CPU_wire_387});
notg #(0, 0) NOT_70 (CPU_wire_388, CPU_wire_86_24);
notg #(0, 0) NOT_71 (CPU_wire_389, CPU_wire_86_25);
notg #(0, 0) NOT_72 (CPU_wire_390, CPU_wire_86_26);
notg #(0, 0) NOT_73 (CPU_wire_391, CPU_wire_86_27);
notg #(0, 0) NOT_74 (CPU_wire_392, CPU_wire_86_28);
notg #(0, 0) NOT_75 (CPU_wire_393, CPU_wire_86_29);
notg #(0, 0) NOT_76 (CPU_wire_394, CPU_wire_86_30);
notg #(0, 0) NOT_77 (CPU_wire_395, CPU_wire_86_31);
and_n #(4, 0, 0) AND_140 (CPU_wire_364, {CPU_wire_86_32, CPU_wire_88_32, CPU_wire_72_0, CPU_wire_8_0});
and_n #(4, 0, 0) AND_141 (CPU_wire_365, {CPU_wire_86_33, CPU_wire_88_33, CPU_wire_70_0, CPU_wire_8_1});
and_n #(4, 0, 0) AND_142 (CPU_wire_366, {CPU_wire_86_34, CPU_wire_88_34, CPU_wire_68_0, CPU_wire_8_2});
and_n #(4, 0, 0) AND_143 (CPU_wire_367, {CPU_wire_86_35, CPU_wire_88_35, CPU_wire_66_0, CPU_wire_8_3});
and_n #(4, 0, 0) AND_144 (CPU_wire_368, {CPU_wire_86_36, CPU_wire_88_36, CPU_wire_64_0, CPU_wire_8_4});
and_n #(4, 0, 0) AND_145 (CPU_wire_369, {CPU_wire_86_37, CPU_wire_88_37, CPU_wire_62_0, CPU_wire_8_5});
and_n #(4, 0, 0) AND_146 (CPU_wire_370, {CPU_wire_86_38, CPU_wire_88_38, CPU_wire_81_0, CPU_wire_8_6});
and_n #(4, 0, 0) AND_147 (CPU_wire_371, {CPU_wire_86_39, CPU_wire_88_39, CPU_wire_80_0, CPU_wire_8_7});
notg #(0, 0) NOT_78 (CPU_wire_396, CPU_wire_86_40);
and_n #(2, 0, 0) AND_148 (CPU_wire_397, {CPU_wire_86_41, CPU_wire_8_8});
notg #(0, 0) NOT_79 (CPU_wire_398, CPU_wire_86_42);
and_n #(3, 0, 0) AND_149 (CPU_wire_399, {CPU_wire_86_43, CPU_wire_88_40, CPU_wire_8_9});
notg #(0, 0) NOT_80 (CPU_wire_373, CPU_wire_88_41);
notg #(0, 0) NOT_81 (CPU_wire_375, CPU_wire_88_42);
notg #(0, 0) NOT_82 (CPU_wire_377, CPU_wire_88_43);
notg #(0, 0) NOT_83 (CPU_wire_379, CPU_wire_88_44);
notg #(0, 0) NOT_84 (CPU_wire_381, CPU_wire_88_45);
notg #(0, 0) NOT_85 (CPU_wire_383, CPU_wire_88_46);
notg #(0, 0) NOT_86 (CPU_wire_385, CPU_wire_88_47);
notg #(0, 0) NOT_87 (CPU_wire_387, CPU_wire_88_48);
and_n #(2, 0, 0) AND_150 (CPU_wire_400, {CPU_wire_88_49, CPU_wire_388});
and_n #(2, 0, 0) AND_151 (CPU_wire_401, {CPU_wire_88_50, CPU_wire_389});
and_n #(2, 0, 0) AND_152 (CPU_wire_402, {CPU_wire_88_51, CPU_wire_390});
and_n #(2, 0, 0) AND_153 (CPU_wire_403, {CPU_wire_88_52, CPU_wire_391});
and_n #(2, 0, 0) AND_154 (CPU_wire_404, {CPU_wire_88_53, CPU_wire_392});
and_n #(2, 0, 0) AND_155 (CPU_wire_405, {CPU_wire_88_54, CPU_wire_393});
and_n #(2, 0, 0) AND_156 (CPU_wire_406, {CPU_wire_88_55, CPU_wire_394});
and_n #(2, 0, 0) AND_157 (CPU_wire_407, {CPU_wire_88_56, CPU_wire_395});
notg #(0, 0) NOT_88 (CPU_wire_408, CPU_wire_88_57);
notg #(0, 0) NOT_89 (CPU_wire_409, CPU_wire_88_58);
and_n #(2, 0, 0) AND_158 (CPU_wire_410, {CPU_wire_88_59, CPU_wire_8_10});
and_n #(2, 0, 0) AND_159 (CPU_wire_411, {CPU_wire_80_1, CPU_wire_8_11});
and_n #(2, 0, 0) AND_160 (CPU_wire_412, {CPU_wire_80_2, CPU_wire_8_12});
and_n #(2, 0, 0) AND_161 (CPU_wire_413, {CPU_wire_80_3, CPU_wire_8_13});
and_n #(2, 0, 0) AND_162 (CPU_wire_414, {CPU_wire_81_1, CPU_wire_8_14});
and_n #(2, 0, 0) AND_163 (CPU_wire_415, {CPU_wire_81_2, CPU_wire_8_15});
and_n #(2, 0, 0) AND_164 (CPU_wire_416, {CPU_wire_81_3, CPU_wire_8_16});
and_n #(2, 0, 0) AND_165 (CPU_wire_417, {CPU_wire_62_1, CPU_wire_8_17});
and_n #(2, 0, 0) AND_166 (CPU_wire_418, {CPU_wire_62_2, CPU_wire_8_18});
and_n #(2, 0, 0) AND_167 (CPU_wire_419, {CPU_wire_62_3, CPU_wire_8_19});
and_n #(2, 0, 0) AND_168 (CPU_wire_420, {CPU_wire_64_1, CPU_wire_8_20});
and_n #(2, 0, 0) AND_169 (CPU_wire_421, {CPU_wire_64_2, CPU_wire_8_21});
and_n #(2, 0, 0) AND_170 (CPU_wire_422, {CPU_wire_64_3, CPU_wire_8_22});
and_n #(2, 0, 0) AND_171 (CPU_wire_423, {CPU_wire_66_1, CPU_wire_8_23});
and_n #(2, 0, 0) AND_172 (CPU_wire_424, {CPU_wire_66_2, CPU_wire_8_24});
and_n #(2, 0, 0) AND_173 (CPU_wire_425, {CPU_wire_66_3, CPU_wire_8_25});
and_n #(2, 0, 0) AND_174 (CPU_wire_426, {CPU_wire_68_1, CPU_wire_8_26});
and_n #(2, 0, 0) AND_175 (CPU_wire_427, {CPU_wire_68_2, CPU_wire_8_27});
and_n #(2, 0, 0) AND_176 (CPU_wire_428, {CPU_wire_68_3, CPU_wire_8_28});
and_n #(2, 0, 0) AND_177 (CPU_wire_429, {CPU_wire_70_1, CPU_wire_8_29});
and_n #(2, 0, 0) AND_178 (CPU_wire_430, {CPU_wire_70_2, CPU_wire_8_30});
and_n #(2, 0, 0) AND_179 (CPU_wire_431, {CPU_wire_70_3, CPU_wire_8_31});
and_n #(2, 0, 0) AND_180 (CPU_wire_432, {CPU_wire_72_1, CPU_wire_8_32});
and_n #(2, 0, 0) AND_181 (CPU_wire_433, {CPU_wire_72_2, CPU_wire_8_33});
and_n #(2, 0, 0) AND_182 (CPU_wire_434, {CPU_wire_72_3, CPU_wire_8_34});
and_n #(3, 0, 0) AND_183 (CPU_wire_435, {CPU_wire_8_35, CPU_wire_396, CPU_wire_408});
and_n #(2, 0, 0) AND_184 (CPU_wire_344, {CPU_wire_411, CPU_wire_436});
nor_n #(2, 0, 0) NOR_1 (CPU_wire_436, {CPU_wire_86_44, CPU_wire_88_60});
and_n #(2, 0, 0) AND_185 (CPU_wire_343, {CPU_wire_414, CPU_wire_437});
nor_n #(2, 0, 0) NOR_2 (CPU_wire_437, {CPU_wire_86_45, CPU_wire_88_61});
and_n #(2, 0, 0) AND_186 (CPU_wire_342, {CPU_wire_417, CPU_wire_438});
nor_n #(2, 0, 0) NOR_3 (CPU_wire_438, {CPU_wire_86_46, CPU_wire_88_62});
and_n #(2, 0, 0) AND_187 (CPU_wire_341, {CPU_wire_420, CPU_wire_439});
nor_n #(2, 0, 0) NOR_4 (CPU_wire_439, {CPU_wire_86_47, CPU_wire_88_63});
and_n #(2, 0, 0) AND_188 (CPU_wire_340, {CPU_wire_423, CPU_wire_440});
nor_n #(2, 0, 0) NOR_5 (CPU_wire_440, {CPU_wire_86_48, CPU_wire_88_64});
and_n #(2, 0, 0) AND_189 (CPU_wire_339, {CPU_wire_426, CPU_wire_441});
nor_n #(2, 0, 0) NOR_6 (CPU_wire_441, {CPU_wire_86_49, CPU_wire_88_65});
and_n #(2, 0, 0) AND_190 (CPU_wire_338, {CPU_wire_429, CPU_wire_442});
nor_n #(2, 0, 0) NOR_7 (CPU_wire_442, {CPU_wire_86_50, CPU_wire_88_66});
and_n #(2, 0, 0) AND_191 (CPU_wire_337, {CPU_wire_432, CPU_wire_443});
nor_n #(2, 0, 0) NOR_8 (CPU_wire_443, {CPU_wire_86_51, CPU_wire_88_67});
or_n #(2, 0, 0) OR_60 (CPU_wire_336, {CPU_wire_435, CPU_wire_110_8});
and_n #(2, 0, 0) AND_192 (CPU_wire_353, {CPU_wire_412, CPU_wire_386});
and_n #(2, 0, 0) AND_193 (CPU_wire_352, {CPU_wire_415, CPU_wire_384});
and_n #(2, 0, 0) AND_194 (CPU_wire_351, {CPU_wire_418, CPU_wire_382});
and_n #(2, 0, 0) AND_195 (CPU_wire_350, {CPU_wire_421, CPU_wire_380});
and_n #(2, 0, 0) AND_196 (CPU_wire_349, {CPU_wire_424, CPU_wire_378});
and_n #(2, 0, 0) AND_197 (CPU_wire_348, {CPU_wire_427, CPU_wire_376});
and_n #(2, 0, 0) AND_198 (CPU_wire_347, {CPU_wire_430, CPU_wire_374});
and_n #(2, 0, 0) AND_199 (CPU_wire_346, {CPU_wire_433, CPU_wire_372});
or_n #(2, 0, 0) OR_61 (CPU_wire_345, {CPU_wire_444, CPU_wire_110_9});
and_n #(2, 0, 0) AND_200 (CPU_wire_444, {CPU_wire_397, CPU_wire_409});
and_n #(2, 0, 0) AND_201 (CPU_wire_362, {CPU_wire_413, CPU_wire_407});
and_n #(2, 0, 0) AND_202 (CPU_wire_361, {CPU_wire_416, CPU_wire_406});
and_n #(2, 0, 0) AND_203 (CPU_wire_360, {CPU_wire_419, CPU_wire_405});
and_n #(2, 0, 0) AND_204 (CPU_wire_359, {CPU_wire_422, CPU_wire_404});
and_n #(2, 0, 0) AND_205 (CPU_wire_358, {CPU_wire_425, CPU_wire_403});
and_n #(2, 0, 0) AND_206 (CPU_wire_357, {CPU_wire_428, CPU_wire_402});
and_n #(2, 0, 0) AND_207 (CPU_wire_356, {CPU_wire_431, CPU_wire_401});
and_n #(2, 0, 0) AND_208 (CPU_wire_355, {CPU_wire_434, CPU_wire_400});
or_n #(2, 0, 0) OR_62 (CPU_wire_354, {CPU_wire_445, CPU_wire_110_10});
and_n #(2, 0, 0) AND_209 (CPU_wire_445, {CPU_wire_410, CPU_wire_398});
or_n #(2, 0, 0) OR_63 (CPU_wire_363, {CPU_wire_399, CPU_wire_110_11});
xor_n #(2, 0, 0) XOR_1 (CPU_wire_446, {CPU_wire_10_1, CPU_wire_12_1});
xor_n #(2, 0, 0) XOR_2 (CPU_wire_447, {CPU_wire_448_0, CPU_wire_14_1});
xor_n #(2, 0, 0) XOR_3 (CPU_wire_449, {CPU_wire_450_0, CPU_wire_16_1});
xor_n #(2, 0, 0) XOR_4 (CPU_wire_451, {CPU_wire_452_0, CPU_wire_18_1});
xor_n #(2, 0, 0) XOR_5 (CPU_wire_453, {CPU_wire_454_0, CPU_wire_20_1});
xor_n #(2, 0, 0) XOR_6 (CPU_wire_455, {CPU_wire_456_0, CPU_wire_22_1});
xor_n #(2, 0, 0) XOR_7 (CPU_wire_457, {CPU_wire_458, CPU_wire_24_1});
and_n #(2, 0, 0) AND_210 (CPU_wire_450, {CPU_wire_448_1, CPU_wire_14_2});
and_n #(2, 0, 0) AND_211 (CPU_wire_448, {CPU_wire_10_2, CPU_wire_12_2});
and_n #(2, 0, 0) AND_212 (CPU_wire_452, {CPU_wire_450_1, CPU_wire_16_2});
and_n #(2, 0, 0) AND_213 (CPU_wire_454, {CPU_wire_452_1, CPU_wire_18_2});
and_n #(2, 0, 0) AND_214 (CPU_wire_456, {CPU_wire_454_1, CPU_wire_20_2});
and_n #(2, 0, 0) AND_215 (CPU_wire_458, {CPU_wire_456_1, CPU_wire_22_2});
and_n #(2, 0, 0) AND_216 (CPU_wire_459, {CPU_wire_6_0, CPU_wire_460});
and_n #(2, 0, 0) AND_217 (CPU_wire_461, {CPU_wire_6_1, CPU_wire_446_0});
and_n #(2, 0, 0) AND_218 (CPU_wire_462, {CPU_wire_6_2, CPU_wire_447_0});
and_n #(2, 0, 0) AND_219 (CPU_wire_463, {CPU_wire_6_3, CPU_wire_449_0});
and_n #(2, 0, 0) AND_220 (CPU_wire_464, {CPU_wire_6_4, CPU_wire_451_0});
and_n #(2, 0, 0) AND_221 (CPU_wire_465, {CPU_wire_6_5, CPU_wire_453_0});
and_n #(2, 0, 0) AND_222 (CPU_wire_466, {CPU_wire_6_6, CPU_wire_455_0});
and_n #(2, 0, 0) AND_223 (CPU_wire_467, {CPU_wire_6_7, CPU_wire_457_0});
and_n #(2, 0, 0) AND_224 (CPU_wire_468, {CPU_wire_6_8, CPU_wire_457_1});
notg #(0, 0) NOT_90 (CPU_wire_469, CPU_wire_6_9);
and_n #(2, 0, 0) AND_225 (CPU_wire_470, {CPU_wire_6_10, CPU_wire_455_1});
notg #(0, 0) NOT_91 (CPU_wire_471, CPU_wire_6_11);
and_n #(2, 0, 0) AND_226 (CPU_wire_472, {CPU_wire_6_12, CPU_wire_453_1});
notg #(0, 0) NOT_92 (CPU_wire_473, CPU_wire_6_13);
and_n #(2, 0, 0) AND_227 (CPU_wire_474, {CPU_wire_6_14, CPU_wire_451_1});
notg #(0, 0) NOT_93 (CPU_wire_475, CPU_wire_6_15);
and_n #(2, 0, 0) AND_228 (CPU_wire_476, {CPU_wire_6_16, CPU_wire_449_1});
notg #(0, 0) NOT_94 (CPU_wire_477, CPU_wire_6_17);
and_n #(2, 0, 0) AND_229 (CPU_wire_478, {CPU_wire_6_18, CPU_wire_447_1});
notg #(0, 0) NOT_95 (CPU_wire_479, CPU_wire_6_19);
and_n #(2, 0, 0) AND_230 (CPU_wire_480, {CPU_wire_6_20, CPU_wire_446_1});
notg #(0, 0) NOT_96 (CPU_wire_481, CPU_wire_6_21);
notg #(0, 0) NOT_97 (CPU_wire_482, CPU_wire_6_22);
and_n #(2, 0, 0) AND_231 (CPU_wire_483, {CPU_wire_6_23, CPU_wire_484});
and_n #(2, 0, 0) AND_232 (CPU_wire_485, {CPU_wire_6_24, CPU_wire_486});
and_n #(2, 0, 0) AND_233 (CPU_wire_487, {CPU_wire_6_25, CPU_wire_10_3});
and_n #(2, 0, 0) AND_234 (CPU_wire_488, {CPU_wire_6_26, CPU_wire_489});
and_n #(2, 0, 0) AND_235 (CPU_wire_490, {CPU_wire_6_27, CPU_wire_491});
and_n #(2, 0, 0) AND_236 (CPU_wire_492, {CPU_wire_6_28, CPU_wire_493});
and_n #(2, 0, 0) AND_237 (CPU_wire_494, {CPU_wire_6_29, CPU_wire_495});
and_n #(2, 0, 0) AND_238 (CPU_wire_496, {CPU_wire_6_30, CPU_wire_497});
and_n #(2, 0, 0) AND_239 (CPU_wire_498, {CPU_wire_6_31, CPU_wire_499});
notg #(0, 0) NOT_98 (CPU_wire_460, CPU_wire_10_4);
notg #(0, 0) NOT_99 (CPU_wire_484, CPU_wire_10_5);
or_n #(2, 0, 0) OR_64 (CPU_wire_500, {CPU_wire_487, CPU_wire_110_12});
or_n #(2, 0, 0) OR_65 (CPU_wire_502, {CPU_wire_485, CPU_wire_110_13});
notg #(0, 0) NOT_100 (CPU_wire_486, CPU_wire_446_2);
or_n #(2, 0, 0) OR_66 (CPU_wire_504, {CPU_wire_488, CPU_wire_110_14});
notg #(0, 0) NOT_101 (CPU_wire_489, CPU_wire_447_2);
or_n #(2, 0, 0) OR_67 (CPU_wire_506, {CPU_wire_490, CPU_wire_110_15});
notg #(0, 0) NOT_102 (CPU_wire_491, CPU_wire_449_2);
or_n #(2, 0, 0) OR_68 (CPU_wire_508, {CPU_wire_492, CPU_wire_110_16});
notg #(0, 0) NOT_103 (CPU_wire_493, CPU_wire_451_2);
or_n #(2, 0, 0) OR_69 (CPU_wire_510, {CPU_wire_494, CPU_wire_110_17});
notg #(0, 0) NOT_104 (CPU_wire_495, CPU_wire_453_2);
or_n #(2, 0, 0) OR_70 (CPU_wire_512, {CPU_wire_496, CPU_wire_110_18});
notg #(0, 0) NOT_105 (CPU_wire_497, CPU_wire_455_2);
or_n #(2, 0, 0) OR_71 (CPU_wire_514, {CPU_wire_498, CPU_wire_110_19});
notg #(0, 0) NOT_106 (CPU_wire_499, CPU_wire_457_2);
or_n #(2, 0, 0) OR_72 (CPU_wire_501, {CPU_wire_516, CPU_wire_483});
and_n #(2, 0, 0) AND_240 (CPU_wire_516, {CPU_wire_482, CPU_wire_49_0});
or_n #(2, 0, 0) OR_73 (CPU_wire_503, {CPU_wire_480, CPU_wire_517});
and_n #(2, 0, 0) AND_241 (CPU_wire_517, {CPU_wire_481, CPU_wire_50_0});
or_n #(2, 0, 0) OR_74 (CPU_wire_505, {CPU_wire_478, CPU_wire_518});
and_n #(2, 0, 0) AND_242 (CPU_wire_518, {CPU_wire_479, CPU_wire_51_0});
or_n #(2, 0, 0) OR_75 (CPU_wire_507, {CPU_wire_476, CPU_wire_519});
and_n #(2, 0, 0) AND_243 (CPU_wire_519, {CPU_wire_477, CPU_wire_52_0});
or_n #(2, 0, 0) OR_76 (CPU_wire_509, {CPU_wire_474, CPU_wire_520});
and_n #(2, 0, 0) AND_244 (CPU_wire_520, {CPU_wire_475, CPU_wire_53_0});
or_n #(2, 0, 0) OR_77 (CPU_wire_511, {CPU_wire_472, CPU_wire_521});
and_n #(2, 0, 0) AND_245 (CPU_wire_521, {CPU_wire_473, CPU_wire_54_0});
or_n #(2, 0, 0) OR_78 (CPU_wire_513, {CPU_wire_470, CPU_wire_522});
and_n #(2, 0, 0) AND_246 (CPU_wire_522, {CPU_wire_471, CPU_wire_55_0});
or_n #(2, 0, 0) OR_79 (CPU_wire_515, {CPU_wire_468, CPU_wire_523});
and_n #(2, 0, 0) AND_247 (CPU_wire_523, {CPU_wire_469, CPU_wire_56_0});
xnor_n #(2, 0, 0) XNOR_1 (CPU_wire_524, {CPU_wire_330_0, CPU_wire_232_0});
xor_n #(2, 0, 0) XOR_8 (CPU_wire_525, {CPU_wire_526, CPU_wire_527});
xnor_n #(2, 0, 0) XNOR_2 (CPU_wire_526, {CPU_wire_120_0, CPU_wire_246_0});
xor_n #(2, 0, 0) XOR_9 (CPU_wire_528, {CPU_wire_529, CPU_wire_530_0});
xnor_n #(2, 0, 0) XNOR_3 (CPU_wire_529, {CPU_wire_136_0, CPU_wire_258_0});
xor_n #(2, 0, 0) XOR_10 (CPU_wire_531, {CPU_wire_532, CPU_wire_533_0});
xnor_n #(2, 0, 0) XNOR_4 (CPU_wire_532, {CPU_wire_152_0, CPU_wire_270_0});
xor_n #(2, 0, 0) XOR_11 (CPU_wire_534, {CPU_wire_535, CPU_wire_536_0});
xnor_n #(2, 0, 0) XNOR_5 (CPU_wire_535, {CPU_wire_168_0, CPU_wire_282_0});
xor_n #(2, 0, 0) XOR_12 (CPU_wire_537, {CPU_wire_538, CPU_wire_539_0});
xnor_n #(2, 0, 0) XNOR_6 (CPU_wire_538, {CPU_wire_184_0, CPU_wire_294_0});
xor_n #(2, 0, 0) XOR_13 (CPU_wire_540, {CPU_wire_541, CPU_wire_542_0});
xnor_n #(2, 0, 0) XNOR_7 (CPU_wire_541, {CPU_wire_200_0, CPU_wire_306_0});
xor_n #(2, 0, 0) XOR_14 (CPU_wire_543, {CPU_wire_544, CPU_wire_545_0});
xnor_n #(2, 0, 0) XNOR_8 (CPU_wire_544, {CPU_wire_216_0, CPU_wire_318_0});
xor_n #(2, 0, 0) XOR_15 (CPU_wire_546, {CPU_wire_330_1, CPU_wire_232_1});
xor_n #(2, 0, 0) XOR_16 (CPU_wire_547, {CPU_wire_548, CPU_wire_549});
xor_n #(2, 0, 0) XOR_17 (CPU_wire_548, {CPU_wire_120_1, CPU_wire_246_1});
xor_n #(2, 0, 0) XOR_18 (CPU_wire_550, {CPU_wire_551, CPU_wire_552_0});
xor_n #(2, 0, 0) XOR_19 (CPU_wire_551, {CPU_wire_136_1, CPU_wire_258_1});
xor_n #(2, 0, 0) XOR_20 (CPU_wire_553, {CPU_wire_554, CPU_wire_555_0});
xor_n #(2, 0, 0) XOR_21 (CPU_wire_554, {CPU_wire_152_1, CPU_wire_270_1});
xor_n #(2, 0, 0) XOR_22 (CPU_wire_556, {CPU_wire_557, CPU_wire_558_0});
xor_n #(2, 0, 0) XOR_23 (CPU_wire_557, {CPU_wire_168_1, CPU_wire_282_1});
xor_n #(2, 0, 0) XOR_24 (CPU_wire_559, {CPU_wire_560, CPU_wire_561_0});
xor_n #(2, 0, 0) XOR_25 (CPU_wire_560, {CPU_wire_184_1, CPU_wire_294_1});
xor_n #(2, 0, 0) XOR_26 (CPU_wire_562, {CPU_wire_563, CPU_wire_564_0});
xor_n #(2, 0, 0) XOR_27 (CPU_wire_563, {CPU_wire_200_1, CPU_wire_306_1});
xor_n #(2, 0, 0) XOR_28 (CPU_wire_565, {CPU_wire_566, CPU_wire_567_0});
xor_n #(2, 0, 0) XOR_29 (CPU_wire_566, {CPU_wire_216_1, CPU_wire_318_1});
and_n #(2, 0, 0) AND_248 (CPU_wire_567, {CPU_wire_232_2, CPU_wire_330_2});
and_n #(2, 0, 0) AND_249 (CPU_wire_568, {CPU_wire_567_1, CPU_wire_318_2});
or_n #(2, 0, 0) OR_80 (CPU_wire_569, {CPU_wire_567_2, CPU_wire_318_3});
or_n #(2, 0, 0) OR_81 (CPU_wire_564, {CPU_wire_568, CPU_wire_570});
and_n #(2, 0, 0) AND_250 (CPU_wire_571, {CPU_wire_564_1, CPU_wire_306_2});
or_n #(2, 0, 0) OR_82 (CPU_wire_572, {CPU_wire_564_2, CPU_wire_306_3});
and_n #(2, 0, 0) AND_251 (CPU_wire_570, {CPU_wire_569, CPU_wire_216_2});
or_n #(2, 0, 0) OR_83 (CPU_wire_561, {CPU_wire_571, CPU_wire_573});
and_n #(2, 0, 0) AND_252 (CPU_wire_574, {CPU_wire_561_1, CPU_wire_294_2});
or_n #(2, 0, 0) OR_84 (CPU_wire_575, {CPU_wire_561_2, CPU_wire_294_3});
and_n #(2, 0, 0) AND_253 (CPU_wire_573, {CPU_wire_572, CPU_wire_200_2});
or_n #(2, 0, 0) OR_85 (CPU_wire_558, {CPU_wire_574, CPU_wire_576});
and_n #(2, 0, 0) AND_254 (CPU_wire_577, {CPU_wire_558_1, CPU_wire_282_2});
or_n #(2, 0, 0) OR_86 (CPU_wire_578, {CPU_wire_558_2, CPU_wire_282_3});
and_n #(2, 0, 0) AND_255 (CPU_wire_576, {CPU_wire_575, CPU_wire_184_2});
or_n #(2, 0, 0) OR_87 (CPU_wire_555, {CPU_wire_577, CPU_wire_579});
and_n #(2, 0, 0) AND_256 (CPU_wire_580, {CPU_wire_555_1, CPU_wire_270_2});
or_n #(2, 0, 0) OR_88 (CPU_wire_581, {CPU_wire_555_2, CPU_wire_270_3});
and_n #(2, 0, 0) AND_257 (CPU_wire_579, {CPU_wire_578, CPU_wire_168_2});
and_n #(2, 0, 0) AND_258 (CPU_wire_582, {CPU_wire_552_1, CPU_wire_258_2});
and_n #(2, 0, 0) AND_259 (CPU_wire_583, {CPU_wire_552_2, CPU_wire_136_2});
or_n #(2, 0, 0) OR_89 (CPU_wire_552, {CPU_wire_580, CPU_wire_584});
and_n #(2, 0, 0) AND_260 (CPU_wire_584, {CPU_wire_581, CPU_wire_152_2});
or_n #(3, 0, 0) OR_90 (CPU_wire_549, {CPU_wire_585, CPU_wire_583, CPU_wire_582});
and_n #(2, 0, 0) AND_261 (CPU_wire_585, {CPU_wire_136_3, CPU_wire_258_3});
or_n #(2, 0, 0) OR_91 (CPU_wire_545, {CPU_wire_586, CPU_wire_232_3});
or_n #(2, 0, 0) OR_92 (CPU_wire_587, {CPU_wire_545_1, CPU_wire_588});
and_n #(2, 0, 0) AND_262 (CPU_wire_589, {CPU_wire_545_2, CPU_wire_590});
notg #(0, 0) NOT_107 (CPU_wire_586, CPU_wire_330_3);
or_n #(2, 0, 0) OR_93 (CPU_wire_542, {CPU_wire_589, CPU_wire_591});
or_n #(2, 0, 0) OR_94 (CPU_wire_592, {CPU_wire_542_1, CPU_wire_593});
and_n #(2, 0, 0) AND_263 (CPU_wire_594, {CPU_wire_542_2, CPU_wire_595});
notg #(0, 0) NOT_108 (CPU_wire_588, CPU_wire_318_4);
notg #(0, 0) NOT_109 (CPU_wire_590, CPU_wire_318_5);
and_n #(2, 0, 0) AND_264 (CPU_wire_591, {CPU_wire_587, CPU_wire_216_3});
or_n #(2, 0, 0) OR_95 (CPU_wire_539, {CPU_wire_594, CPU_wire_596});
or_n #(2, 0, 0) OR_96 (CPU_wire_597, {CPU_wire_539_1, CPU_wire_598});
and_n #(2, 0, 0) AND_265 (CPU_wire_599, {CPU_wire_539_2, CPU_wire_600});
notg #(0, 0) NOT_110 (CPU_wire_593, CPU_wire_306_4);
notg #(0, 0) NOT_111 (CPU_wire_595, CPU_wire_306_5);
and_n #(2, 0, 0) AND_266 (CPU_wire_596, {CPU_wire_592, CPU_wire_200_3});
or_n #(2, 0, 0) OR_97 (CPU_wire_536, {CPU_wire_599, CPU_wire_601});
or_n #(2, 0, 0) OR_98 (CPU_wire_602, {CPU_wire_536_1, CPU_wire_603});
and_n #(2, 0, 0) AND_267 (CPU_wire_604, {CPU_wire_536_2, CPU_wire_605});
notg #(0, 0) NOT_112 (CPU_wire_598, CPU_wire_294_4);
notg #(0, 0) NOT_113 (CPU_wire_600, CPU_wire_294_5);
and_n #(2, 0, 0) AND_268 (CPU_wire_601, {CPU_wire_597, CPU_wire_184_3});
or_n #(2, 0, 0) OR_99 (CPU_wire_533, {CPU_wire_604, CPU_wire_606});
or_n #(2, 0, 0) OR_100 (CPU_wire_607, {CPU_wire_533_1, CPU_wire_608});
and_n #(2, 0, 0) AND_269 (CPU_wire_609, {CPU_wire_533_2, CPU_wire_610});
notg #(0, 0) NOT_114 (CPU_wire_603, CPU_wire_282_4);
notg #(0, 0) NOT_115 (CPU_wire_605, CPU_wire_282_5);
and_n #(2, 0, 0) AND_270 (CPU_wire_606, {CPU_wire_602, CPU_wire_168_3});
and_n #(2, 0, 0) AND_271 (CPU_wire_611, {CPU_wire_530_1, CPU_wire_612});
and_n #(2, 0, 0) AND_272 (CPU_wire_613, {CPU_wire_530_2, CPU_wire_136_4});
or_n #(2, 0, 0) OR_101 (CPU_wire_530, {CPU_wire_609, CPU_wire_614});
notg #(0, 0) NOT_116 (CPU_wire_608, CPU_wire_270_4);
notg #(0, 0) NOT_117 (CPU_wire_610, CPU_wire_270_5);
and_n #(2, 0, 0) AND_273 (CPU_wire_614, {CPU_wire_607, CPU_wire_152_3});
or_n #(3, 0, 0) OR_102 (CPU_wire_527, {CPU_wire_615, CPU_wire_613, CPU_wire_611});
and_n #(2, 0, 0) AND_274 (CPU_wire_615, {CPU_wire_616, CPU_wire_136_5});
notg #(0, 0) NOT_118 (CPU_wire_616, CPU_wire_258_4);
notg #(0, 0) NOT_119 (CPU_wire_612, CPU_wire_258_5);
nor_n #(2, 0, 0) NOR_9 (CPU_wire_617, {CPU_wire_2_1, CPU_wire_4_2});
and_n #(2, 0, 0) AND_275 (CPU_wire_620, {CPU_wire_619_0, CPU_wire_642_0});
or_n #(2, 0, 0) OR_103 (CPU_wire_618, {CPU_wire_643, CPU_wire_644});
and_n #(2, 0, 0) AND_276 (CPU_wire_643, {CPU_wire_2_2, CPU_wire_4_3});
notg #(0, 0) NOT_120 (CPU_wire_645, CPU_wire_619_1);
and_n #(2, 0, 0) AND_277 (CPU_wire_644, {CPU_wire_645, CPU_wire_642_1});
and_n #(2, 0, 0) AND_278 (CPU_wire_623, {CPU_wire_622_0, CPU_wire_642_2});
or_n #(2, 0, 0) OR_104 (CPU_wire_621, {CPU_wire_646, CPU_wire_647});
and_n #(2, 0, 0) AND_279 (CPU_wire_646, {CPU_wire_2_3, CPU_wire_4_4});
notg #(0, 0) NOT_121 (CPU_wire_648, CPU_wire_622_1);
and_n #(2, 0, 0) AND_280 (CPU_wire_647, {CPU_wire_648, CPU_wire_642_3});
and_n #(2, 0, 0) AND_281 (CPU_wire_626, {CPU_wire_625_0, CPU_wire_642_4});
or_n #(2, 0, 0) OR_105 (CPU_wire_624, {CPU_wire_649, CPU_wire_650});
and_n #(2, 0, 0) AND_282 (CPU_wire_649, {CPU_wire_2_4, CPU_wire_4_5});
notg #(0, 0) NOT_122 (CPU_wire_651, CPU_wire_625_1);
and_n #(2, 0, 0) AND_283 (CPU_wire_650, {CPU_wire_651, CPU_wire_642_5});
and_n #(2, 0, 0) AND_284 (CPU_wire_629, {CPU_wire_628_0, CPU_wire_642_6});
or_n #(2, 0, 0) OR_106 (CPU_wire_627, {CPU_wire_652, CPU_wire_653});
and_n #(2, 0, 0) AND_285 (CPU_wire_652, {CPU_wire_2_5, CPU_wire_4_6});
notg #(0, 0) NOT_123 (CPU_wire_654, CPU_wire_628_1);
and_n #(2, 0, 0) AND_286 (CPU_wire_653, {CPU_wire_654, CPU_wire_642_7});
and_n #(2, 0, 0) AND_287 (CPU_wire_632, {CPU_wire_631_0, CPU_wire_642_8});
or_n #(2, 0, 0) OR_107 (CPU_wire_630, {CPU_wire_655, CPU_wire_656});
and_n #(2, 0, 0) AND_288 (CPU_wire_655, {CPU_wire_2_6, CPU_wire_4_7});
notg #(0, 0) NOT_124 (CPU_wire_657, CPU_wire_631_1);
and_n #(2, 0, 0) AND_289 (CPU_wire_656, {CPU_wire_657, CPU_wire_642_9});
and_n #(2, 0, 0) AND_290 (CPU_wire_635, {CPU_wire_634_0, CPU_wire_642_10});
or_n #(2, 0, 0) OR_108 (CPU_wire_633, {CPU_wire_658, CPU_wire_659});
and_n #(2, 0, 0) AND_291 (CPU_wire_658, {CPU_wire_2_7, CPU_wire_4_8});
notg #(0, 0) NOT_125 (CPU_wire_660, CPU_wire_634_1);
and_n #(2, 0, 0) AND_292 (CPU_wire_659, {CPU_wire_660, CPU_wire_642_11});
and_n #(2, 0, 0) AND_293 (CPU_wire_638, {CPU_wire_637_0, CPU_wire_642_12});
or_n #(2, 0, 0) OR_109 (CPU_wire_636, {CPU_wire_661, CPU_wire_662});
and_n #(2, 0, 0) AND_294 (CPU_wire_661, {CPU_wire_2_8, CPU_wire_4_9});
notg #(0, 0) NOT_126 (CPU_wire_663, CPU_wire_637_1);
and_n #(2, 0, 0) AND_295 (CPU_wire_662, {CPU_wire_663, CPU_wire_642_13});
and_n #(2, 0, 0) AND_296 (CPU_wire_641, {CPU_wire_640_0, CPU_wire_642_14});
or_n #(2, 0, 0) OR_110 (CPU_wire_639, {CPU_wire_664, CPU_wire_665});
and_n #(2, 0, 0) AND_297 (CPU_wire_664, {CPU_wire_2_9, CPU_wire_4_10});
notg #(0, 0) NOT_127 (CPU_wire_666, CPU_wire_640_1);
and_n #(2, 0, 0) AND_298 (CPU_wire_665, {CPU_wire_666, CPU_wire_642_15});
and_n #(2, 0, 0) AND_299 (CPU_wire_667, {CPU_wire_546, CPU_wire_668});
and_n #(2, 0, 0) AND_300 (CPU_wire_669, {CPU_wire_565, CPU_wire_670});
and_n #(2, 0, 0) AND_301 (CPU_wire_671, {CPU_wire_562, CPU_wire_672});
and_n #(2, 0, 0) AND_302 (CPU_wire_673, {CPU_wire_559, CPU_wire_674});
and_n #(2, 0, 0) AND_303 (CPU_wire_675, {CPU_wire_556, CPU_wire_676});
and_n #(2, 0, 0) AND_304 (CPU_wire_677, {CPU_wire_553, CPU_wire_678});
and_n #(2, 0, 0) AND_305 (CPU_wire_679, {CPU_wire_550, CPU_wire_680});
and_n #(2, 0, 0) AND_306 (CPU_wire_681, {CPU_wire_547, CPU_wire_682});
or_n #(2, 0, 0) OR_111 (CPU_wire_619, {CPU_wire_667, CPU_wire_683});
and_n #(2, 0, 0) AND_307 (CPU_wire_684, {CPU_wire_232_4, CPU_wire_685_0});
or_n #(2, 0, 0) OR_112 (CPU_wire_686, {CPU_wire_684, CPU_wire_687});
nor_n #(2, 0, 0) NOR_10 (CPU_wire_687, {CPU_wire_524, CPU_wire_685_1});
notg #(0, 0) NOT_128 (CPU_wire_668, CPU_wire_642_16);
and_n #(2, 0, 0) AND_308 (CPU_wire_683, {CPU_wire_686, CPU_wire_642_17});
or_n #(2, 0, 0) OR_113 (CPU_wire_622, {CPU_wire_669, CPU_wire_688});
and_n #(2, 0, 0) AND_309 (CPU_wire_689, {CPU_wire_216_4, CPU_wire_685_2});
or_n #(2, 0, 0) OR_114 (CPU_wire_690, {CPU_wire_689, CPU_wire_691});
notg #(0, 0) NOT_129 (CPU_wire_692, CPU_wire_685_3);
and_n #(2, 0, 0) AND_310 (CPU_wire_691, {CPU_wire_692, CPU_wire_543});
notg #(0, 0) NOT_130 (CPU_wire_670, CPU_wire_642_18);
and_n #(2, 0, 0) AND_311 (CPU_wire_688, {CPU_wire_690, CPU_wire_642_19});
or_n #(2, 0, 0) OR_115 (CPU_wire_625, {CPU_wire_671, CPU_wire_693});
and_n #(2, 0, 0) AND_312 (CPU_wire_694, {CPU_wire_200_4, CPU_wire_685_4});
or_n #(2, 0, 0) OR_116 (CPU_wire_695, {CPU_wire_694, CPU_wire_696});
notg #(0, 0) NOT_131 (CPU_wire_697, CPU_wire_685_5);
and_n #(2, 0, 0) AND_313 (CPU_wire_696, {CPU_wire_697, CPU_wire_540});
notg #(0, 0) NOT_132 (CPU_wire_672, CPU_wire_642_20);
and_n #(2, 0, 0) AND_314 (CPU_wire_693, {CPU_wire_695, CPU_wire_642_21});
or_n #(2, 0, 0) OR_117 (CPU_wire_628, {CPU_wire_673, CPU_wire_698});
and_n #(2, 0, 0) AND_315 (CPU_wire_699, {CPU_wire_184_4, CPU_wire_685_6});
or_n #(2, 0, 0) OR_118 (CPU_wire_700, {CPU_wire_699, CPU_wire_701});
notg #(0, 0) NOT_133 (CPU_wire_702, CPU_wire_685_7);
and_n #(2, 0, 0) AND_316 (CPU_wire_701, {CPU_wire_702, CPU_wire_537});
notg #(0, 0) NOT_134 (CPU_wire_674, CPU_wire_642_22);
and_n #(2, 0, 0) AND_317 (CPU_wire_698, {CPU_wire_700, CPU_wire_642_23});
or_n #(2, 0, 0) OR_119 (CPU_wire_631, {CPU_wire_675, CPU_wire_703});
and_n #(2, 0, 0) AND_318 (CPU_wire_704, {CPU_wire_168_4, CPU_wire_685_8});
or_n #(2, 0, 0) OR_120 (CPU_wire_705, {CPU_wire_704, CPU_wire_706});
notg #(0, 0) NOT_135 (CPU_wire_707, CPU_wire_685_9);
and_n #(2, 0, 0) AND_319 (CPU_wire_706, {CPU_wire_707, CPU_wire_534});
notg #(0, 0) NOT_136 (CPU_wire_676, CPU_wire_642_24);
and_n #(2, 0, 0) AND_320 (CPU_wire_703, {CPU_wire_705, CPU_wire_642_25});
or_n #(2, 0, 0) OR_121 (CPU_wire_634, {CPU_wire_677, CPU_wire_708});
and_n #(2, 0, 0) AND_321 (CPU_wire_709, {CPU_wire_152_4, CPU_wire_685_10});
or_n #(2, 0, 0) OR_122 (CPU_wire_710, {CPU_wire_709, CPU_wire_711});
notg #(0, 0) NOT_137 (CPU_wire_712, CPU_wire_685_11);
and_n #(2, 0, 0) AND_322 (CPU_wire_711, {CPU_wire_712, CPU_wire_531});
notg #(0, 0) NOT_138 (CPU_wire_678, CPU_wire_642_26);
and_n #(2, 0, 0) AND_323 (CPU_wire_708, {CPU_wire_710, CPU_wire_642_27});
or_n #(2, 0, 0) OR_123 (CPU_wire_637, {CPU_wire_679, CPU_wire_713});
and_n #(2, 0, 0) AND_324 (CPU_wire_714, {CPU_wire_136_6, CPU_wire_685_12});
or_n #(2, 0, 0) OR_124 (CPU_wire_715, {CPU_wire_714, CPU_wire_716});
notg #(0, 0) NOT_139 (CPU_wire_717, CPU_wire_685_13);
and_n #(2, 0, 0) AND_325 (CPU_wire_716, {CPU_wire_717, CPU_wire_528});
notg #(0, 0) NOT_140 (CPU_wire_680, CPU_wire_642_28);
and_n #(2, 0, 0) AND_326 (CPU_wire_713, {CPU_wire_715, CPU_wire_642_29});
or_n #(2, 0, 0) OR_125 (CPU_wire_640, {CPU_wire_681, CPU_wire_718});
and_n #(2, 0, 0) AND_327 (CPU_wire_719, {CPU_wire_120_2, CPU_wire_685_14});
or_n #(2, 0, 0) OR_126 (CPU_wire_720, {CPU_wire_719, CPU_wire_721});
notg #(0, 0) NOT_141 (CPU_wire_722, CPU_wire_685_15);
and_n #(2, 0, 0) AND_328 (CPU_wire_721, {CPU_wire_722, CPU_wire_525});
notg #(0, 0) NOT_142 (CPU_wire_682, CPU_wire_642_30);
and_n #(2, 0, 0) AND_329 (CPU_wire_718, {CPU_wire_720, CPU_wire_642_31});
xor_n #(2, 0, 0) XOR_30 (CPU_wire_642, {CPU_wire_2_10, CPU_wire_4_11});
notg #(0, 0) NOT_143 (CPU_wire_723, CPU_wire_2_11);
and_n #(2, 0, 0) AND_330 (CPU_wire_685, {CPU_wire_4_12, CPU_wire_723});
xor_n #(2, 0, 0) XOR_31 (CPU_wire_26, {CPU_wire_75_17, CPU_wire_10_6});
xor_n #(2, 0, 0) XOR_32 (CPU_wire_47, {CPU_wire_724, CPU_wire_725});
xor_n #(2, 0, 0) XOR_33 (CPU_wire_44, {CPU_wire_726, CPU_wire_727_0});
xor_n #(2, 0, 0) XOR_34 (CPU_wire_41, {CPU_wire_728, CPU_wire_729_0});
xor_n #(2, 0, 0) XOR_35 (CPU_wire_38, {CPU_wire_730, CPU_wire_731_0});
xor_n #(2, 0, 0) XOR_36 (CPU_wire_35, {CPU_wire_732, CPU_wire_733_0});
xor_n #(2, 0, 0) XOR_37 (CPU_wire_732, {CPU_wire_16_3, CPU_wire_88_68});
xor_n #(2, 0, 0) XOR_38 (CPU_wire_32, {CPU_wire_734, CPU_wire_735_0});
xor_n #(2, 0, 0) XOR_39 (CPU_wire_734, {CPU_wire_14_3, CPU_wire_86_52});
xor_n #(2, 0, 0) XOR_40 (CPU_wire_29, {CPU_wire_736, CPU_wire_737_0});
xor_n #(2, 0, 0) XOR_41 (CPU_wire_736, {CPU_wire_12_3, CPU_wire_78_33});
bufg #(0, 0) BUF_2 (CPU_wire_730, CPU_wire_18_3);
bufg #(0, 0) BUF_3 (CPU_wire_728, CPU_wire_20_3);
bufg #(0, 0) BUF_4 (CPU_wire_726, CPU_wire_22_3);
bufg #(0, 0) BUF_5 (CPU_wire_724, CPU_wire_24_2);
and_n #(2, 0, 0) AND_331 (CPU_wire_737, {CPU_wire_10_7, CPU_wire_75_18});
and_n #(2, 0, 0) AND_332 (CPU_wire_738, {CPU_wire_737_1, CPU_wire_78_34});
or_n #(2, 0, 0) OR_127 (CPU_wire_739, {CPU_wire_737_2, CPU_wire_78_35});
or_n #(2, 0, 0) OR_128 (CPU_wire_735, {CPU_wire_738, CPU_wire_740});
and_n #(2, 0, 0) AND_333 (CPU_wire_741, {CPU_wire_735_1, CPU_wire_86_53});
or_n #(2, 0, 0) OR_129 (CPU_wire_742, {CPU_wire_735_2, CPU_wire_86_54});
and_n #(2, 0, 0) AND_334 (CPU_wire_740, {CPU_wire_739, CPU_wire_12_4});
or_n #(2, 0, 0) OR_130 (CPU_wire_733, {CPU_wire_741, CPU_wire_743});
and_n #(2, 0, 0) AND_335 (CPU_wire_744, {CPU_wire_733_1, CPU_wire_88_69});
or_n #(2, 0, 0) OR_131 (CPU_wire_745, {CPU_wire_733_2, CPU_wire_88_70});
and_n #(2, 0, 0) AND_336 (CPU_wire_743, {CPU_wire_742, CPU_wire_14_4});
or_n #(2, 0, 0) OR_132 (CPU_wire_731, {CPU_wire_744, CPU_wire_746});
and_n #(2, 0, 0) AND_337 (CPU_wire_729, {CPU_wire_731_1, CPU_wire_18_4});
and_n #(2, 0, 0) AND_338 (CPU_wire_746, {CPU_wire_745, CPU_wire_16_4});
and_n #(2, 0, 0) AND_339 (CPU_wire_727, {CPU_wire_729_1, CPU_wire_20_4});
and_n #(2, 0, 0) AND_340 (CPU_wire_725, {CPU_wire_727_1, CPU_wire_22_4});
bufg #(0, 0) BUF_6 (address_7, CPU_wire_49_1);
bufg #(0, 0) BUF_7 (address_6, CPU_wire_50_1);
bufg #(0, 0) BUF_8 (address_5, CPU_wire_51_1);
bufg #(0, 0) BUF_9 (address_4, CPU_wire_52_1);
bufg #(0, 0) BUF_10 (address_3, CPU_wire_53_1);
bufg #(0, 0) BUF_11 (address_2, CPU_wire_54_1);
bufg #(0, 0) BUF_12 (address_1, CPU_wire_55_1);
bufg #(0, 0) BUF_13 (address_0, CPU_wire_56_1);
bufg #(0, 0) BUF_14 (CPU_wire_82, clk_net_0);
bufg #(0, 0) BUF_15 (CPU_wire_94, inst_7);
bufg #(0, 0) BUF_16 (CPU_wire_96, inst_6);
bufg #(0, 0) BUF_17 (CPU_wire_98, inst_5);
bufg #(0, 0) BUF_18 (CPU_wire_100, inst_4);
bufg #(0, 0) BUF_19 (CPU_wire_102, inst_3);
bufg #(0, 0) BUF_20 (CPU_wire_104, inst_2);
bufg #(0, 0) BUF_21 (CPU_wire_106, inst_1);
bufg #(0, 0) BUF_22 (CPU_wire_108, inst_0);
bufg #(0, 0) BUF_23 (out_data_7, CPU_wire_58_1);
bufg #(0, 0) BUF_24 (out_data_6, CPU_wire_61_1);
bufg #(0, 0) BUF_25 (out_data_5, CPU_wire_63_1);
bufg #(0, 0) BUF_26 (out_data_4, CPU_wire_65_1);
bufg #(0, 0) BUF_27 (out_data_3, CPU_wire_67_1);
bufg #(0, 0) BUF_28 (out_data_2, CPU_wire_69_1);
bufg #(0, 0) BUF_29 (out_data_1, CPU_wire_71_1);
bufg #(0, 0) BUF_30 (out_data_0, CPU_wire_73_1);
bufg #(0, 0) BUF_31 (CPU_wire_110, reset_net_0);
bufg #(0, 0) BUF_32 (store_net_0, CPU_wire_3);

/*
dff DFF_1  (CPU_wire_75, CPU_wire_83, CPU_wire_82, 1'b0, 1'b0, 1'b1, NbarT, Si, 1'b0);
dff DFF_2  (CPU_wire_78, CPU_wire_84, CPU_wire_82, 1'b0, 1'b0, 1'b1, NbarT, Si, 1'b0);
dff DFF_3  (CPU_wire_86, CPU_wire_85, CPU_wire_82, 1'b0, 1'b0, 1'b1, NbarT, Si, 1'b0);
dff DFF_4  (CPU_wire_88, CPU_wire_87, CPU_wire_82, 1'b0, 1'b0, 1'b1, NbarT, Si, 1'b0);
dff DFF_5  (CPU_wire_2, CPU_wire_89, CPU_wire_82, 1'b0, 1'b0, 1'b1, NbarT, Si, 1'b0);
dff DFF_6  (CPU_wire_4, CPU_wire_90, CPU_wire_82, 1'b0, 1'b0, 1'b1, NbarT, Si, 1'b0);
dff DFF_7  (CPU_wire_92, CPU_wire_91, CPU_wire_82, 1'b0, 1'b0, 1'b1, NbarT, Si, 1'b0);
dff DFF_8  (CPU_wire_7, CPU_wire_93, CPU_wire_82, 1'b0, 1'b0, 1'b1, NbarT, Si, 1'b0);
dff DFF_9  (CPU_wire_126, CPU_wire_337, CPU_wire_82, CPU_wire_335, 1'b0, CPU_wire_336, NbarT, Si, 1'b0);
dff DFF_10  (CPU_wire_142, CPU_wire_338, CPU_wire_82, CPU_wire_335, 1'b0, CPU_wire_336, NbarT, Si, 1'b0);
dff DFF_11  (CPU_wire_158, CPU_wire_339, CPU_wire_82, CPU_wire_335, 1'b0, CPU_wire_336, NbarT, Si, 1'b0);
dff DFF_12  (CPU_wire_174, CPU_wire_340, CPU_wire_82, CPU_wire_335, 1'b0, CPU_wire_336, NbarT, Si, 1'b0);
dff DFF_13  (CPU_wire_190, CPU_wire_341, CPU_wire_82, CPU_wire_335, 1'b0, CPU_wire_336, NbarT, Si, 1'b0);
dff DFF_14  (CPU_wire_206, CPU_wire_342, CPU_wire_82, CPU_wire_335, 1'b0, CPU_wire_336, NbarT, Si, 1'b0);
dff DFF_15  (CPU_wire_222, CPU_wire_343, CPU_wire_82, CPU_wire_335, 1'b0, CPU_wire_336, NbarT, Si, 1'b0);
dff DFF_16  (CPU_wire_238, CPU_wire_344, CPU_wire_82, CPU_wire_335, 1'b0, CPU_wire_336, NbarT, Si, 1'b0);
dff DFF_17  (CPU_wire_116, CPU_wire_346, CPU_wire_82, CPU_wire_335, 1'b0, CPU_wire_345, NbarT, Si, 1'b0);
dff DFF_18  (CPU_wire_132, CPU_wire_347, CPU_wire_82, CPU_wire_335, 1'b0, CPU_wire_345, NbarT, Si, 1'b0);
dff DFF_19  (CPU_wire_148, CPU_wire_348, CPU_wire_82, CPU_wire_335, 1'b0, CPU_wire_345, NbarT, Si, 1'b0);
dff DFF_20  (CPU_wire_164, CPU_wire_349, CPU_wire_82, CPU_wire_335, 1'b0, CPU_wire_345, NbarT, Si, 1'b0);
dff DFF_21  (CPU_wire_180, CPU_wire_350, CPU_wire_82, CPU_wire_335, 1'b0, CPU_wire_345, NbarT, Si, 1'b0);
dff DFF_22  (CPU_wire_196, CPU_wire_351, CPU_wire_82, CPU_wire_335, 1'b0, CPU_wire_345, NbarT, Si, 1'b0);
dff DFF_23  (CPU_wire_212, CPU_wire_352, CPU_wire_82, CPU_wire_335, 1'b0, CPU_wire_345, NbarT, Si, 1'b0);
dff DFF_24  (CPU_wire_228, CPU_wire_353, CPU_wire_82, CPU_wire_335, 1'b0, CPU_wire_345, NbarT, Si, 1'b0);
dff DFF_25  (CPU_wire_123, CPU_wire_355, CPU_wire_82, CPU_wire_335, 1'b0, CPU_wire_354, NbarT, Si, 1'b0);
dff DFF_26  (CPU_wire_139, CPU_wire_356, CPU_wire_82, CPU_wire_335, 1'b0, CPU_wire_354, NbarT, Si, 1'b0);
dff DFF_27  (CPU_wire_155, CPU_wire_357, CPU_wire_82, CPU_wire_335, 1'b0, CPU_wire_354, NbarT, Si, 1'b0);
dff DFF_28  (CPU_wire_171, CPU_wire_358, CPU_wire_82, CPU_wire_335, 1'b0, CPU_wire_354, NbarT, Si, 1'b0);
dff DFF_29  (CPU_wire_187, CPU_wire_359, CPU_wire_82, CPU_wire_335, 1'b0, CPU_wire_354, NbarT, Si, 1'b0);
dff DFF_30  (CPU_wire_203, CPU_wire_360, CPU_wire_82, CPU_wire_335, 1'b0, CPU_wire_354, NbarT, Si, 1'b0);
dff DFF_31  (CPU_wire_219, CPU_wire_361, CPU_wire_82, CPU_wire_335, 1'b0, CPU_wire_354, NbarT, Si, 1'b0);
dff DFF_32  (CPU_wire_235, CPU_wire_362, CPU_wire_82, CPU_wire_335, 1'b0, CPU_wire_354, NbarT, Si, 1'b0);
dff DFF_33  (CPU_wire_112, CPU_wire_364, CPU_wire_82, CPU_wire_335, 1'b0, CPU_wire_363, NbarT, Si, 1'b0);
dff DFF_34  (CPU_wire_128, CPU_wire_365, CPU_wire_82, CPU_wire_335, 1'b0, CPU_wire_363, NbarT, Si, 1'b0);
dff DFF_35  (CPU_wire_144, CPU_wire_366, CPU_wire_82, CPU_wire_335, 1'b0, CPU_wire_363, NbarT, Si, 1'b0);
dff DFF_36  (CPU_wire_160, CPU_wire_367, CPU_wire_82, CPU_wire_335, 1'b0, CPU_wire_363, NbarT, Si, 1'b0);
dff DFF_37  (CPU_wire_176, CPU_wire_368, CPU_wire_82, CPU_wire_335, 1'b0, CPU_wire_363, NbarT, Si, 1'b0);
dff DFF_38  (CPU_wire_192, CPU_wire_369, CPU_wire_82, CPU_wire_335, 1'b0, CPU_wire_363, NbarT, Si, 1'b0);
dff DFF_39  (CPU_wire_208, CPU_wire_370, CPU_wire_82, CPU_wire_335, 1'b0, CPU_wire_363, NbarT, Si, 1'b0);
dff DFF_40  (CPU_wire_224, CPU_wire_371, CPU_wire_82, CPU_wire_335, 1'b0, CPU_wire_363, NbarT, Si, 1'b0);
dff DFF_41  (CPU_wire_10, CPU_wire_501, CPU_wire_7, CPU_wire_500, CPU_wire_459, CE, NbarT, Si, 1'b0);
dff DFF_42  (CPU_wire_12, CPU_wire_503, CPU_wire_7, CPU_wire_502, CPU_wire_461, CE, NbarT, Si, 1'b0);
dff DFF_43  (CPU_wire_14, CPU_wire_505, CPU_wire_7, CPU_wire_504, CPU_wire_462, CE, NbarT, Si, 1'b0);
dff DFF_44  (CPU_wire_16, CPU_wire_507, CPU_wire_7, CPU_wire_506, CPU_wire_463, CE, NbarT, Si, 1'b0);
dff DFF_45  (CPU_wire_18, CPU_wire_509, CPU_wire_7, CPU_wire_508, CPU_wire_464, CE, NbarT, Si, 1'b0);
dff DFF_46  (CPU_wire_20, CPU_wire_511, CPU_wire_7, CPU_wire_510, CPU_wire_465, CE, NbarT, Si, 1'b0);
dff DFF_47  (CPU_wire_22, CPU_wire_513, CPU_wire_7, CPU_wire_512, CPU_wire_466, CE, NbarT, Si, 1'b0);
dff DFF_48  (CPU_wire_24, CPU_wire_515, CPU_wire_7, CPU_wire_514, CPU_wire_467, CE, NbarT, Si, 1'b0);
dff DFF_49  (CPU_wire_58, CPU_wire_619, CPU_wire_617, CPU_wire_618, CPU_wire_620, CE, NbarT, Si, 1'b0);
dff DFF_50  (CPU_wire_61, CPU_wire_622, CPU_wire_617, CPU_wire_621, CPU_wire_623, CE, NbarT, Si, 1'b0);
dff DFF_51  (CPU_wire_63, CPU_wire_625, CPU_wire_617, CPU_wire_624, CPU_wire_626, CE, NbarT, Si, 1'b0);
dff DFF_52  (CPU_wire_65, CPU_wire_628, CPU_wire_617, CPU_wire_627, CPU_wire_629, CE, NbarT, Si, 1'b0);
dff DFF_53  (CPU_wire_67, CPU_wire_631, CPU_wire_617, CPU_wire_630, CPU_wire_632, CE, NbarT, Si, 1'b0);
dff DFF_54  (CPU_wire_69, CPU_wire_634, CPU_wire_617, CPU_wire_633, CPU_wire_635, CE, NbarT, Si, 1'b0);
dff DFF_55  (CPU_wire_71, CPU_wire_637, CPU_wire_617, CPU_wire_636, CPU_wire_638, CE, NbarT, Si, 1'b0);
dff DFF_56  (CPU_wire_73, CPU_wire_640, CPU_wire_617, CPU_wire_639, CPU_wire_641, CE, NbarT, Si, 1'b0);
*/
endmodule
